* SPICE NETLIST
***************************************

.SUBCKT n12ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT p12ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT n18ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT p18ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT nt12ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT nt18ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT nhvt12ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT phvt12ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT nlvt12LL_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT plvt12ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT n12ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT n12ll_ckt_rf_sdc DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT n18ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT nlvt12ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT nlvt12ll_ckt_rf_sdc DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw12ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw12ll_ckt_rf_sdc DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnwlvt12ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnwlvt12ll_ckt_rf_sdc DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw18ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p12ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p12ll_ckt_rf_sdc DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT plvt12ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT plvt12ll_ckt_rf_sdc DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p18ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT n12ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT n12ll_ckt_rf_sdc_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT nlvt12ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT nlvt12ll_ckt_rf_sdc_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p12ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p12ll_ckt_rf_sdc_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT plvt12ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT plvt12ll_ckt_rf_sdc_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw12ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw12ll_ckt_rf_sdc_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnwlvt12ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnwlvt12ll_ckt_rf_sdc_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT n18ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p18ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw18ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw12ll_ckt D G S B
.ENDS
***************************************
.SUBCKT dnw18ll_ckt D G S B
.ENDS
***************************************
.SUBCKT dnwhvt12ll_ckt D G S B
.ENDS
***************************************
.SUBCKT dnwlvt12ll_ckt D G S B
.ENDS
***************************************
.SUBCKT n25ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT p25ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT nt25ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT ntod33ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT nod33ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT pod33ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT n25ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT n25llod33_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT n25llod33_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT n25ll_ckt_rf_sdc DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT n25ll_ckt_rf_sdc_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw25ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw25llod33_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw25llod33_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw25ll_ckt_rf_sdc DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw25ll_ckt_rf_sdc_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p25ll_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p25llod33_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p25llod33_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p25ll_ckt_rf_sdc DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p25ll_ckt_rf_sdc_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw25ll_ckt D G S B
.ENDS
***************************************
.SUBCKT dnwod33ll_ckt D G S B
.ENDS
***************************************
.SUBCKT dnwud18ll_ckt D G S B
.ENDS
***************************************
.SUBCKT n25ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT p25ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw25ll_ckt_rf_mis DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT pvar12ll_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar12ll_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar12ll_ckt_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT pvar12lldnw_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar12lldnw_ckt_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT pvar18ll_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar18ll_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar18ll_ckt_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT pvar18lldnw_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar18lldnw_ckt_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT pvardio12ll_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvardio18ll_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar25ll_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar25ll_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar25ll_ckt_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT pvar25lldnw_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar25lldnw_ckt_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT pvardio25ll_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT rndifsab_ckt_rf PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpdifsab_ckt_rf PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnposab_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT rnposab_ckt_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpposab_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT rpposab_ckt_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT rndif_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpdif_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT rppo_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwsti_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwaa_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rndifsab_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpdifsab_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnposab_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT rpposab_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpo_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnposab_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpposab_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rm1_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rm2_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rm3_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rm4_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT ralpa_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rm5_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rm6_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rtm1_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT rtm2_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom13_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT mom13_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom13_wops_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom24_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT mom24_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom24_wops_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom14_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT mom14_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom14_wops_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom15_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT mom15_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom15_wops_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom25_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT mom25_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom25_wops_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom35_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT mom35_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom35_wops_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom16_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT mom16_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom16_wops_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom26_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT mom26_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom26_wops_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom36_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT mom36_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom36_wops_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom46_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT mom46_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom46_wops_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mom13_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom14_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom24_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom15_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom25_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom35_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom16_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom26_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom36_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom46_3t_ckt PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom13_wops_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom24_wops_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom14_wops_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom15_wops_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom25_wops_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom35_wops_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom16_wops_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom26_wops_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom36_wops_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom46_wops_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom13_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom24_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom14_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom15_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom25_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom35_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom16_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom26_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom36_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT mom46_rf_3t PLUS MINUS B
.ENDS
***************************************
.SUBCKT nld50ll_ckt D G S B
.ENDS
***************************************
.SUBCKT pld50ll_ckt D G S B
.ENDS
***************************************
.SUBCKT nld50ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT pld50ll_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT nld50llod_ckt D G S B
.ENDS
***************************************
.SUBCKT pld50llod_ckt D G S B
.ENDS
***************************************
.SUBCKT nld50llod_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT pld50llod_mis_ckt D G S B
.ENDS
***************************************
.SUBCKT 65smic_062swl_svt_strap_v0p0
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT 65smic_062swl_svt_edge_v0p0 1 2 3 6 7 8
** N=8 EP=6 IP=0 FDC=3
M0 7 1 3 1 DNNPGSVT L=7.5e-08 W=1.25e-07 $X=965 $Y=90 $D=96
M1 6 1 1 1 DNNPDSVT L=6.5e-08 W=2.1e-07 $X=125 $Y=90 $D=95
M2 8 1 2 2 DNPLSVT L=6.5e-08 W=9.5e-08 $X=470 $Y=90 $D=97
.ENDS
***************************************
.SUBCKT 65smic_062swl_svt_dummycell_v0p0 1 2 3 4 5
** N=11 EP=5 IP=0 FDC=6
M0 3 1 8 2 DNNPGSVT L=7.5e-08 W=1.25e-07 $X=150 $Y=335 $D=96
M1 9 2 5 2 DNNPGSVT L=7.5e-08 W=1.25e-07 $X=965 $Y=90 $D=96
M2 8 9 2 2 DNNPDSVT L=6.5e-08 W=2.1e-07 $X=125 $Y=90 $D=95
M3 2 8 9 2 DNNPDSVT L=6.5e-08 W=2.1e-07 $X=905 $Y=345 $D=95
M4 8 9 4 4 DNPLSVT L=6.5e-08 W=9.5e-08 $X=470 $Y=90 $D=97
M5 4 8 9 4 DNPLSVT L=6.5e-08 W=9.5e-08 $X=675 $Y=345 $D=97
.ENDS
***************************************
.SUBCKT bitcell_dummy_lr_2B_620_VHSSP 1 2 3 4 5 6
** N=9 EP=6 IP=14 FDC=12
X0 1 2 3 4 9 65smic_062swl_svt_dummycell_v0p0 $T=0 500 1 0 $X=-125 $Y=-185
X1 5 2 6 4 9 65smic_062swl_svt_dummycell_v0p0 $T=0 500 0 0 $X=-125 $Y=315
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6 7 8
** N=11 EP=8 IP=16 FDC=24
X0 2 1 4 5 3 11 bitcell_dummy_lr_2B_620_VHSSP $T=0 0 0 0 $X=-125 $Y=-185
X1 6 1 11 5 7 8 bitcell_dummy_lr_2B_620_VHSSP $T=0 1000 0 0 $X=-125 $Y=815
.ENDS
***************************************
.SUBCKT bitcell_dummy_lr_2A_620_VHSSP 1 2 3 4 5 6
** N=9 EP=6 IP=14 FDC=12
X0 1 2 9 3 4 65smic_062swl_svt_dummycell_v0p0 $T=0 0 0 0 $X=-125 $Y=-185
X1 5 2 9 3 6 65smic_062swl_svt_dummycell_v0p0 $T=0 1000 1 0 $X=-125 $Y=315
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8
** N=11 EP=8 IP=16 FDC=24
X0 1 3 4 5 2 11 bitcell_dummy_lr_2A_620_VHSSP $T=0 0 0 0 $X=-125 $Y=-185
X1 6 3 4 11 7 8 bitcell_dummy_lr_2A_620_VHSSP $T=0 1000 0 0 $X=-125 $Y=815
.ENDS
***************************************
.SUBCKT bitcell64_dummy_620_VHSSP 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67
** N=100 EP=67 IP=212 FDC=408
X3 1 2 68 89 95 97 65smic_062swl_svt_edge_v0p0 $T=0 950 1 0 $X=-125 $Y=394
X4 1 2 69 90 96 98 65smic_062swl_svt_edge_v0p0 $T=0 17950 0 0 $X=-125 $Y=17765
X5 1 2 70 93 91 99 65smic_062swl_svt_edge_v0p0 $T=1240 19150 0 180 $X=-125 $Y=18594
X6 1 2 71 94 92 100 65smic_062swl_svt_edge_v0p0 $T=1240 35150 1 180 $X=-125 $Y=34965
X7 1 3 4 70 2 5 6 72 ICV_1 $T=0 19150 0 0 $X=-125 $Y=18965
X8 1 7 8 72 2 9 10 73 ICV_1 $T=0 21150 0 0 $X=-125 $Y=20965
X9 1 11 12 73 2 13 14 74 ICV_1 $T=0 23150 0 0 $X=-125 $Y=22965
X10 1 15 16 74 2 17 18 75 ICV_1 $T=0 25150 0 0 $X=-125 $Y=24965
X11 1 19 20 75 2 21 22 76 ICV_1 $T=0 27150 0 0 $X=-125 $Y=26965
X12 1 23 24 76 2 25 26 77 ICV_1 $T=0 29150 0 0 $X=-125 $Y=28965
X13 1 27 28 77 2 29 30 78 ICV_1 $T=0 31150 0 0 $X=-125 $Y=30965
X14 1 31 32 78 2 33 34 71 ICV_1 $T=0 33150 0 0 $X=-125 $Y=32965
X15 35 1 2 79 36 69 bitcell_dummy_lr_2A_620_VHSSP $T=0 16950 0 0 $X=-125 $Y=16765
X16 1 37 1 2 68 38 39 80 ICV_2 $T=0 950 0 0 $X=-125 $Y=765
X17 40 41 1 2 80 42 43 81 ICV_2 $T=0 2950 0 0 $X=-125 $Y=2765
X18 44 45 1 2 81 46 47 82 ICV_2 $T=0 4950 0 0 $X=-125 $Y=4765
X19 48 49 1 2 82 50 51 83 ICV_2 $T=0 6950 0 0 $X=-125 $Y=6765
X20 52 53 1 2 83 54 55 84 ICV_2 $T=0 8950 0 0 $X=-125 $Y=8765
X21 56 57 1 2 84 58 59 85 ICV_2 $T=0 10950 0 0 $X=-125 $Y=10765
X22 60 61 1 2 85 62 63 86 ICV_2 $T=0 12950 0 0 $X=-125 $Y=12765
X23 64 65 1 2 86 66 67 79 ICV_2 $T=0 14950 0 0 $X=-125 $Y=14765
.ENDS
***************************************
.SUBCKT YMUX8_CAP_LEFT_620
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT Y8_DOWN_POWER_BW_620
** N=37 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD DATA DOUT BWEN
.ENDS
***************************************
.SUBCKT smic_062_strap_x2_VHSSP
** N=6 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT smic_062_edge_x2b_VHSSP 1 2 3 4 7 8 9 10 11 12
** N=12 EP=10 IP=16 FDC=6
X0 1 2 3 7 8 11 65smic_062swl_svt_edge_v0p0 $T=1240 0 1 180 $X=-125 $Y=-185
X1 1 2 4 9 10 12 65smic_062swl_svt_edge_v0p0 $T=1240 0 0 0 $X=1115 $Y=-185
.ENDS
***************************************
.SUBCKT 65smic_062swl_svt_bitcell_v0p0 1 2 3 4 5
** N=9 EP=5 IP=0 FDC=6
M0 3 1 6 2 DNNPGSVT L=7.5e-08 W=1.25e-07 $X=150 $Y=335 $D=96
M1 7 1 5 2 DNNPGSVT L=7.5e-08 W=1.25e-07 $X=965 $Y=90 $D=96
M2 6 7 2 2 DNNPDSVT L=6.5e-08 W=2.1e-07 $X=125 $Y=90 $D=95
M3 2 6 7 2 DNNPDSVT L=6.5e-08 W=2.1e-07 $X=905 $Y=345 $D=95
M4 6 7 4 4 DNPLSVT L=6.5e-08 W=9.5e-08 $X=470 $Y=90 $D=97
M5 4 6 7 4 DNPLSVT L=6.5e-08 W=9.5e-08 $X=675 $Y=345 $D=97
.ENDS
***************************************
.SUBCKT smic_062_bitcellx4b_VHSSP 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=20 FDC=24
X0 1 2 3 4 5 65smic_062swl_svt_bitcell_v0p0 $T=1240 0 1 180 $X=-125 $Y=-185
X1 6 2 3 4 5 65smic_062swl_svt_bitcell_v0p0 $T=1240 1000 0 180 $X=-125 $Y=315
X2 1 2 7 4 8 65smic_062swl_svt_bitcell_v0p0 $T=1240 0 0 0 $X=1115 $Y=-185
X3 6 2 7 4 8 65smic_062swl_svt_bitcell_v0p0 $T=1240 1000 1 0 $X=1115 $Y=315
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=16 FDC=48
X0 2 1 9 5 4 3 10 6 smic_062_bitcellx4b_VHSSP $T=0 0 0 0 $X=-125 $Y=-185
X1 7 1 9 5 4 8 10 6 smic_062_bitcellx4b_VHSSP $T=0 1000 0 0 $X=-125 $Y=815
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7 8 9 10 11 12 13 14
** N=14 EP=14 IP=20 FDC=96
X0 1 2 3 6 7 8 4 5 13 14 ICV_3 $T=0 0 0 0 $X=-125 $Y=-185
X1 1 9 10 6 7 8 11 12 13 14 ICV_3 $T=0 2000 0 0 $X=-125 $Y=1815
.ENDS
***************************************
.SUBCKT smic_062_edge_x2a_VHSSP 1 2 3 4 7 8 9 10 11 12
** N=12 EP=10 IP=16 FDC=6
X0 1 2 3 7 8 11 65smic_062swl_svt_edge_v0p0 $T=0 0 0 0 $X=-125 $Y=-185
X1 1 2 4 9 10 12 65smic_062swl_svt_edge_v0p0 $T=2480 0 1 180 $X=1115 $Y=-185
.ENDS
***************************************
.SUBCKT smic_062_bitcellx4a_VHSSP 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=20 FDC=24
X0 1 2 3 4 5 65smic_062swl_svt_bitcell_v0p0 $T=0 0 0 0 $X=-125 $Y=-185
X1 6 2 3 4 5 65smic_062swl_svt_bitcell_v0p0 $T=0 1000 1 0 $X=-125 $Y=315
X2 1 2 7 4 8 65smic_062swl_svt_bitcell_v0p0 $T=2480 0 1 180 $X=1115 $Y=-185
X3 6 2 7 4 8 65smic_062swl_svt_bitcell_v0p0 $T=2480 1000 0 180 $X=1115 $Y=315
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=16 FDC=48
X0 1 3 9 4 5 2 10 6 smic_062_bitcellx4a_VHSSP $T=0 0 0 0 $X=-125 $Y=-185
X1 7 3 9 4 5 8 10 6 smic_062_bitcellx4a_VHSSP $T=0 1000 0 0 $X=-125 $Y=815
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8 9 10 11 12 13 14
** N=14 EP=14 IP=20 FDC=96
X0 2 3 1 6 7 8 4 5 13 14 ICV_5 $T=0 0 0 0 $X=-125 $Y=-185
X1 9 10 1 6 7 8 11 12 13 14 ICV_5 $T=0 2000 0 0 $X=-125 $Y=1815
.ENDS
***************************************
.SUBCKT a_x64y2_ab_620_VHSSP 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71
** N=95 EP=71 IP=186 FDC=816
X3 1 3 2 4 76 74 80 86 90 92 smic_062_edge_x2b_VHSSP $T=0 19150 1 0 $X=-125 $Y=18594
X4 1 3 2 4 77 75 81 87 91 93 smic_062_edge_x2b_VHSSP $T=0 35150 0 0 $X=-125 $Y=34965
X5 1 5 6 7 8 2 3 4 9 10 11 12 37 38 ICV_4 $T=0 19150 0 0 $X=-125 $Y=18965
X6 1 13 14 15 16 2 3 4 17 18 19 20 37 38 ICV_4 $T=0 23150 0 0 $X=-125 $Y=22965
X7 1 21 22 23 24 2 3 4 25 26 27 28 37 38 ICV_4 $T=0 27150 0 0 $X=-125 $Y=26965
X8 1 29 30 31 32 2 3 4 33 34 35 36 37 38 ICV_4 $T=0 31150 0 0 $X=-125 $Y=30965
X9 1 3 37 38 72 78 84 82 88 94 smic_062_edge_x2a_VHSSP $T=0 950 1 0 $X=-125 $Y=394
X10 1 3 37 38 73 79 85 83 89 95 smic_062_edge_x2a_VHSSP $T=0 17950 0 0 $X=-125 $Y=17765
X11 39 1 2 3 37 40 4 38 smic_062_bitcellx4a_VHSSP $T=0 16950 0 0 $X=-125 $Y=16765
X12 1 1 41 42 43 3 37 38 44 45 46 47 2 4 ICV_6 $T=0 950 0 0 $X=-125 $Y=765
X13 1 48 49 50 51 3 37 38 52 53 54 55 2 4 ICV_6 $T=0 4950 0 0 $X=-125 $Y=4765
X14 1 56 57 58 59 3 37 38 60 61 62 63 2 4 ICV_6 $T=0 8950 0 0 $X=-125 $Y=8765
X15 1 64 65 66 67 3 37 38 68 69 70 71 2 4 ICV_6 $T=0 12950 0 0 $X=-125 $Y=12765
.ENDS
***************************************
.SUBCKT Y8_X64_1_DOWN_BW_620_VHSSP 1 2 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43
+ 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85
** N=85 EP=82 IP=289 FDC=3264
X1 1 70 2 73 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53
+ 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 71 72 36 37
+ 1 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35
+ a_x64y2_ab_620_VHSSP $T=0 0 0 0 $X=-125 $Y=-285
X2 1 74 2 77 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53
+ 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 75 76 36 37
+ 1 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35
+ a_x64y2_ab_620_VHSSP $T=2480 0 0 0 $X=2355 $Y=-285
X3 1 78 2 81 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53
+ 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 79 80 36 37
+ 1 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35
+ a_x64y2_ab_620_VHSSP $T=4960 0 0 0 $X=4835 $Y=-285
X4 1 82 2 85 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53
+ 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 83 84 36 37
+ 1 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35
+ a_x64y2_ab_620_VHSSP $T=7440 0 0 0 $X=7315 $Y=-285
.ENDS
***************************************
.SUBCKT Y8_TOP_POWER_620
** N=34 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT Y8_X64_1_UP_620_VHSSP 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83
** N=86 EP=83 IP=286 FDC=3264
X0 1 68 67 71 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 69 70 33 34
+ 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32
+ a_x64y2_ab_620_VHSSP $T=0 0 0 0 $X=-125 $Y=-285
X1 1 72 67 75 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 73 74 33 34
+ 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32
+ a_x64y2_ab_620_VHSSP $T=2480 0 0 0 $X=2355 $Y=-285
X2 1 76 67 79 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 77 78 33 34
+ 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32
+ a_x64y2_ab_620_VHSSP $T=4960 0 0 0 $X=4835 $Y=-285
X3 1 80 67 83 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 81 82 33 34
+ 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32
+ a_x64y2_ab_620_VHSSP $T=7440 0 0 0 $X=7315 $Y=-285
.ENDS
***************************************
.SUBCKT YMX8SAWR_BW_620 VSS VDD LBL[0] UBL[0] LBLX[0] UBLX[0] YX[1] YX[0] DATA LBLX[1] UBLX[1] LBL[1] UBL[1] YX[2] LBL[2] UBL[2] WE LBLX[2] UBLX[2] CLK
+ CLKX LBLX[3] UBLX[3] LBL[3] UBL[3] YX[3] YX[5] DOUT LBL[4] UBL[4] AXS LBLX[4] UBLX[4] AS LBLX[5] UBLX[5] LBL[5] UBL[5] LBL[6] UBL[6]
+ YX[6] LBLX[6] UBLX[6] SACK1 YX[4] LBLX[7] UBLX[7] LBL[7] UBL[7] SACK4 BWEN YX[7]
** N=227 EP=52 IP=0 FDC=377
M0 LBL[0] 95 61 VSS n12ll L=6e-08 W=7.5e-07 $X=395 $Y=2800 $D=0
M1 61 95 LBL[0] VSS n12ll L=6e-08 W=7.5e-07 $X=395 $Y=3080 $D=0
M2 LBLX[0] 72 61 VSS n12ll L=6e-08 W=7.5e-07 $X=395 $Y=3360 $D=0
M3 61 72 LBLX[0] VSS n12ll L=6e-08 W=7.5e-07 $X=395 $Y=3640 $D=0
M4 UBLX[0] 72 62 VSS n12ll L=6e-08 W=7.5e-07 $X=395 $Y=29670 $D=0
M5 62 72 UBLX[0] VSS n12ll L=6e-08 W=7.5e-07 $X=395 $Y=29950 $D=0
M6 UBL[0] 95 62 VSS n12ll L=6e-08 W=7.5e-07 $X=395 $Y=30230 $D=0
M7 62 95 UBL[0] VSS n12ll L=6e-08 W=7.5e-07 $X=395 $Y=30510 $D=0
M8 VSS 63 57 VSS n12ll L=6e-08 W=8e-07 $X=445 $Y=5385 $D=0
M9 VSS 64 58 VSS n12ll L=6e-08 W=8e-07 $X=445 $Y=27185 $D=0
M10 VSS 57 61 VSS n12ll L=6e-08 W=1.52e-06 $X=490 $Y=4590 $D=0
M11 68 74 VSS VSS n12ll L=6e-08 W=1.52e-06 $X=490 $Y=4860 $D=0
M12 VSS 75 69 VSS n12ll L=6e-08 W=1.52e-06 $X=490 $Y=28450 $D=0
M13 62 58 VSS VSS n12ll L=6e-08 W=1.52e-06 $X=490 $Y=28720 $D=0
M14 185 60 VSS VSS n12ll L=6e-08 W=8e-07 $X=725 $Y=5385 $D=0
M15 186 60 VSS VSS n12ll L=6e-08 W=8e-07 $X=725 $Y=27185 $D=0
M16 63 65 185 VSS n12ll L=6e-08 W=8e-07 $X=925 $Y=5385 $D=0
M17 64 66 186 VSS n12ll L=6e-08 W=8e-07 $X=925 $Y=27185 $D=0
M18 LBL[1] 95 68 VSS n12ll L=6e-08 W=7.5e-07 $X=1335 $Y=2800 $D=0
M19 68 95 LBL[1] VSS n12ll L=6e-08 W=7.5e-07 $X=1335 $Y=3080 $D=0
M20 LBLX[1] 72 68 VSS n12ll L=6e-08 W=7.5e-07 $X=1335 $Y=3360 $D=0
M21 68 72 LBLX[1] VSS n12ll L=6e-08 W=7.5e-07 $X=1335 $Y=3640 $D=0
M22 UBLX[1] 72 69 VSS n12ll L=6e-08 W=7.5e-07 $X=1335 $Y=29670 $D=0
M23 69 72 UBLX[1] VSS n12ll L=6e-08 W=7.5e-07 $X=1335 $Y=29950 $D=0
M24 UBL[1] 95 69 VSS n12ll L=6e-08 W=7.5e-07 $X=1335 $Y=30230 $D=0
M25 69 95 UBL[1] VSS n12ll L=6e-08 W=7.5e-07 $X=1335 $Y=30510 $D=0
M26 VSS VSS DATA VSS n12ll L=6e-08 W=2e-07 $X=1410 $Y=16190 $D=0
M27 VSS DATA 67 VSS n12ll L=6e-08 W=4e-07 $X=1445 $Y=12440 $D=0
M28 187 65 70 VSS n12ll L=6e-08 W=8e-07 $X=1495 $Y=5385 $D=0
M29 188 66 71 VSS n12ll L=6e-08 W=8e-07 $X=1495 $Y=27185 $D=0
M30 VSS YX[0] 60 VSS n12ll L=6e-08 W=4e-07 $X=1675 $Y=22905 $D=0
M31 59 YX[1] VSS VSS n12ll L=6e-08 W=4e-07 $X=1685 $Y=10365 $D=0
M32 VSS 59 187 VSS n12ll L=6e-08 W=8e-07 $X=1695 $Y=5385 $D=0
M33 VSS 59 188 VSS n12ll L=6e-08 W=8e-07 $X=1695 $Y=27185 $D=0
M34 72 77 VSS VSS n12ll L=6e-08 W=1e-06 $X=1790 $Y=18090 $D=0
M35 76 67 VSS VSS n12ll L=3e-07 W=4e-07 $X=1835 $Y=12440 $D=0
M36 73 91 VSS VSS n12ll L=6e-08 W=4e-07 $X=1860 $Y=16110 $D=0
M37 74 70 VSS VSS n12ll L=6e-08 W=8e-07 $X=1975 $Y=5385 $D=0
M38 75 71 VSS VSS n12ll L=6e-08 W=8e-07 $X=1975 $Y=27185 $D=0
M39 VSS 77 72 VSS n12ll L=6e-08 W=1e-06 $X=2080 $Y=18090 $D=0
M40 189 73 VSS VSS n12ll L=6e-08 W=1e-06 $X=2415 $Y=18090 $D=0
M41 VSS 83 80 VSS n12ll L=6e-08 W=5e-07 $X=2510 $Y=16135 $D=0
M42 77 80 189 VSS n12ll L=6e-08 W=1e-06 $X=2635 $Y=18090 $D=0
M43 190 WE VSS VSS n12ll L=6e-08 W=4e-07 $X=2800 $Y=16135 $D=0
M44 VSS 76 84 VSS n12ll L=2e-07 W=4e-07 $X=2845 $Y=12440 $D=0
M45 LBL[2] 95 85 VSS n12ll L=6e-08 W=7.5e-07 $X=2875 $Y=2800 $D=0
M46 85 95 LBL[2] VSS n12ll L=6e-08 W=7.5e-07 $X=2875 $Y=3080 $D=0
M47 LBLX[2] 72 85 VSS n12ll L=6e-08 W=7.5e-07 $X=2875 $Y=3360 $D=0
M48 85 72 LBLX[2] VSS n12ll L=6e-08 W=7.5e-07 $X=2875 $Y=3640 $D=0
M49 UBLX[2] 72 86 VSS n12ll L=6e-08 W=7.5e-07 $X=2875 $Y=29670 $D=0
M50 86 72 UBLX[2] VSS n12ll L=6e-08 W=7.5e-07 $X=2875 $Y=29950 $D=0
M51 UBL[2] 95 86 VSS n12ll L=6e-08 W=7.5e-07 $X=2875 $Y=30230 $D=0
M52 86 95 UBL[2] VSS n12ll L=6e-08 W=7.5e-07 $X=2875 $Y=30510 $D=0
M53 VSS 87 78 VSS n12ll L=6e-08 W=8e-07 $X=2925 $Y=5385 $D=0
M54 VSS 88 79 VSS n12ll L=6e-08 W=8e-07 $X=2925 $Y=27185 $D=0
M55 VSS YX[2] 82 VSS n12ll L=6e-08 W=4e-07 $X=2960 $Y=10455 $D=0
M56 81 YX[3] VSS VSS n12ll L=6e-08 W=4e-07 $X=2960 $Y=10745 $D=0
M57 VSS 78 85 VSS n12ll L=6e-08 W=1.52e-06 $X=2970 $Y=4590 $D=0
M58 92 98 VSS VSS n12ll L=6e-08 W=1.52e-06 $X=2970 $Y=4860 $D=0
M59 VSS 99 93 VSS n12ll L=6e-08 W=1.52e-06 $X=2970 $Y=28450 $D=0
M60 86 79 VSS VSS n12ll L=6e-08 W=1.52e-06 $X=2970 $Y=28720 $D=0
M61 83 101 190 VSS n12ll L=6e-08 W=4e-07 $X=3030 $Y=16135 $D=0
M62 191 82 VSS VSS n12ll L=6e-08 W=8e-07 $X=3205 $Y=5385 $D=0
M63 192 82 VSS VSS n12ll L=6e-08 W=8e-07 $X=3205 $Y=27185 $D=0
M64 193 80 90 VSS n12ll L=6e-08 W=1e-06 $X=3255 $Y=18090 $D=0
M65 89 84 VSS VSS n12ll L=6e-08 W=7e-07 $X=3355 $Y=12195 $D=0
M66 87 65 191 VSS n12ll L=6e-08 W=8e-07 $X=3405 $Y=5385 $D=0
M67 88 66 192 VSS n12ll L=6e-08 W=8e-07 $X=3405 $Y=27185 $D=0
M68 VSS 91 193 VSS n12ll L=6e-08 W=1e-06 $X=3475 $Y=18090 $D=0
M69 94 CLKX 89 VSS n12ll L=6e-08 W=7e-07 $X=3700 $Y=12195 $D=0
M70 95 90 VSS VSS n12ll L=6e-08 W=1e-06 $X=3805 $Y=18090 $D=0
M71 LBL[3] 95 92 VSS n12ll L=6e-08 W=7.5e-07 $X=3815 $Y=2800 $D=0
M72 92 95 LBL[3] VSS n12ll L=6e-08 W=7.5e-07 $X=3815 $Y=3080 $D=0
M73 LBLX[3] 72 92 VSS n12ll L=6e-08 W=7.5e-07 $X=3815 $Y=3360 $D=0
M74 92 72 LBLX[3] VSS n12ll L=6e-08 W=7.5e-07 $X=3815 $Y=3640 $D=0
M75 UBLX[3] 72 93 VSS n12ll L=6e-08 W=7.5e-07 $X=3815 $Y=29670 $D=0
M76 93 72 UBLX[3] VSS n12ll L=6e-08 W=7.5e-07 $X=3815 $Y=29950 $D=0
M77 UBL[3] 95 93 VSS n12ll L=6e-08 W=7.5e-07 $X=3815 $Y=30230 $D=0
M78 93 95 UBL[3] VSS n12ll L=6e-08 W=7.5e-07 $X=3815 $Y=30510 $D=0
M79 194 65 96 VSS n12ll L=6e-08 W=8e-07 $X=3975 $Y=5385 $D=0
M80 195 66 97 VSS n12ll L=6e-08 W=8e-07 $X=3975 $Y=27185 $D=0
M81 VSS 91 94 VSS n12ll L=6e-07 W=1.2e-07 $X=4075 $Y=11570 $D=0
M82 VSS 90 95 VSS n12ll L=6e-08 W=1e-06 $X=4095 $Y=18090 $D=0
M83 VSS 81 194 VSS n12ll L=6e-08 W=8e-07 $X=4175 $Y=5385 $D=0
M84 VSS 81 195 VSS n12ll L=6e-08 W=8e-07 $X=4175 $Y=27185 $D=0
M85 98 96 VSS VSS n12ll L=6e-08 W=8e-07 $X=4455 $Y=5385 $D=0
M86 99 97 VSS VSS n12ll L=6e-08 W=8e-07 $X=4455 $Y=27185 $D=0
M87 VSS 94 91 VSS n12ll L=6e-08 W=5e-07 $X=4485 $Y=12205 $D=0
M88 VSS 109 DOUT VSS n12ll L=6e-08 W=5e-07 $X=4675 $Y=16425 $D=0
M89 DOUT 109 VSS VSS n12ll L=6e-08 W=5e-07 $X=4965 $Y=16425 $D=0
M90 110 101 VSS VSS n12ll L=6e-07 W=1.2e-07 $X=5045 $Y=11625 $D=0
M91 VSS 109 DOUT VSS n12ll L=6e-08 W=5e-07 $X=5255 $Y=16425 $D=0
M92 VSS AXS 66 VSS n12ll L=6e-08 W=4e-07 $X=5305 $Y=22645 $D=0
M93 102 YX[5] VSS VSS n12ll L=6e-08 W=4e-07 $X=5305 $Y=22990 $D=0
M94 VSS 110 101 VSS n12ll L=6e-08 W=4e-07 $X=5345 $Y=12275 $D=0
M95 LBL[4] 95 106 VSS n12ll L=6e-08 W=7.5e-07 $X=5355 $Y=2800 $D=0
M96 106 95 LBL[4] VSS n12ll L=6e-08 W=7.5e-07 $X=5355 $Y=3080 $D=0
M97 LBLX[4] 72 106 VSS n12ll L=6e-08 W=7.5e-07 $X=5355 $Y=3360 $D=0
M98 106 72 LBLX[4] VSS n12ll L=6e-08 W=7.5e-07 $X=5355 $Y=3640 $D=0
M99 UBLX[4] 72 107 VSS n12ll L=6e-08 W=7.5e-07 $X=5355 $Y=29670 $D=0
M100 107 72 UBLX[4] VSS n12ll L=6e-08 W=7.5e-07 $X=5355 $Y=29950 $D=0
M101 UBL[4] 95 107 VSS n12ll L=6e-08 W=7.5e-07 $X=5355 $Y=30230 $D=0
M102 107 95 UBL[4] VSS n12ll L=6e-08 W=7.5e-07 $X=5355 $Y=30510 $D=0
M103 VSS 111 103 VSS n12ll L=6e-08 W=8e-07 $X=5405 $Y=5385 $D=0
M104 VSS 112 104 VSS n12ll L=6e-08 W=8e-07 $X=5405 $Y=27185 $D=0
M105 VSS 103 106 VSS n12ll L=6e-08 W=1.52e-06 $X=5450 $Y=4590 $D=0
M106 115 123 VSS VSS n12ll L=6e-08 W=1.52e-06 $X=5450 $Y=4860 $D=0
M107 VSS 124 116 VSS n12ll L=6e-08 W=1.52e-06 $X=5450 $Y=28450 $D=0
M108 107 104 VSS VSS n12ll L=6e-08 W=1.52e-06 $X=5450 $Y=28720 $D=0
M109 108 100 125 VSS n12ll L=1e-07 W=1.5e-06 $X=5460 $Y=17605 $D=0
M110 196 100 VSS VSS n12ll L=6e-08 W=1e-06 $X=5595 $Y=16050 $D=0
M111 197 105 VSS VSS n12ll L=6e-08 W=8e-07 $X=5685 $Y=5385 $D=0
M112 198 105 VSS VSS n12ll L=6e-08 W=8e-07 $X=5685 $Y=27185 $D=0
M113 109 119 196 VSS n12ll L=6e-08 W=1e-06 $X=5835 $Y=16050 $D=0
M114 111 65 197 VSS n12ll L=6e-08 W=8e-07 $X=5885 $Y=5385 $D=0
M115 112 66 198 VSS n12ll L=6e-08 W=8e-07 $X=5885 $Y=27185 $D=0
M116 125 100 108 VSS n12ll L=1e-07 W=1.5e-06 $X=5920 $Y=17605 $D=0
M117 114 CLKX 110 VSS n12ll L=6e-08 W=7e-07 $X=6120 $Y=12140 $D=0
M118 LBL[5] 95 115 VSS n12ll L=6e-08 W=7.5e-07 $X=6295 $Y=2800 $D=0
M119 115 95 LBL[5] VSS n12ll L=6e-08 W=7.5e-07 $X=6295 $Y=3080 $D=0
M120 LBLX[5] 72 115 VSS n12ll L=6e-08 W=7.5e-07 $X=6295 $Y=3360 $D=0
M121 115 72 LBLX[5] VSS n12ll L=6e-08 W=7.5e-07 $X=6295 $Y=3640 $D=0
M122 UBLX[5] 72 116 VSS n12ll L=6e-08 W=7.5e-07 $X=6295 $Y=29670 $D=0
M123 116 72 UBLX[5] VSS n12ll L=6e-08 W=7.5e-07 $X=6295 $Y=29950 $D=0
M124 UBL[5] 95 116 VSS n12ll L=6e-08 W=7.5e-07 $X=6295 $Y=30230 $D=0
M125 116 95 UBL[5] VSS n12ll L=6e-08 W=7.5e-07 $X=6295 $Y=30510 $D=0
M126 100 108 125 VSS n12ll L=1e-07 W=1.5e-06 $X=6380 $Y=17605 $D=0
M127 199 65 117 VSS n12ll L=6e-08 W=8e-07 $X=6455 $Y=5385 $D=0
M128 200 66 118 VSS n12ll L=6e-08 W=8e-07 $X=6455 $Y=27185 $D=0
M129 VSS 122 114 VSS n12ll L=6e-08 W=7e-07 $X=6490 $Y=12140 $D=0
M130 201 109 119 VSS n12ll L=6e-08 W=1e-06 $X=6515 $Y=16050 $D=0
M131 VSS YX[4] 105 VSS n12ll L=6e-08 W=3.95e-07 $X=6585 $Y=10330 $D=0
M132 65 AS VSS VSS n12ll L=6e-08 W=3.95e-07 $X=6585 $Y=10630 $D=0
M133 VSS 102 199 VSS n12ll L=6e-08 W=8e-07 $X=6655 $Y=5385 $D=0
M134 VSS 102 200 VSS n12ll L=6e-08 W=8e-07 $X=6655 $Y=27185 $D=0
M135 VSS 108 201 VSS n12ll L=6e-08 W=1e-06 $X=6805 $Y=16050 $D=0
M136 122 127 VSS VSS n12ll L=2e-07 W=4e-07 $X=6830 $Y=12440 $D=0
M137 125 108 100 VSS n12ll L=1e-07 W=1.5e-06 $X=6840 $Y=17605 $D=0
M138 123 117 VSS VSS n12ll L=6e-08 W=8e-07 $X=6935 $Y=5385 $D=0
M139 124 118 VSS VSS n12ll L=6e-08 W=8e-07 $X=6935 $Y=27185 $D=0
M140 VSS 130 126 VSS n12ll L=6e-08 W=5e-07 $X=7465 $Y=16135 $D=0
M141 VSS 135 127 VSS n12ll L=3e-07 W=4e-07 $X=7735 $Y=12440 $D=0
M142 130 SACK1 VSS VSS n12ll L=6e-08 W=4e-07 $X=7755 $Y=16135 $D=0
M143 LBL[6] 95 133 VSS n12ll L=6e-08 W=7.5e-07 $X=7835 $Y=2800 $D=0
M144 133 95 LBL[6] VSS n12ll L=6e-08 W=7.5e-07 $X=7835 $Y=3080 $D=0
M145 LBLX[6] 72 133 VSS n12ll L=6e-08 W=7.5e-07 $X=7835 $Y=3360 $D=0
M146 133 72 LBLX[6] VSS n12ll L=6e-08 W=7.5e-07 $X=7835 $Y=3640 $D=0
M147 UBLX[6] 72 134 VSS n12ll L=6e-08 W=7.5e-07 $X=7835 $Y=29670 $D=0
M148 134 72 UBLX[6] VSS n12ll L=6e-08 W=7.5e-07 $X=7835 $Y=29950 $D=0
M149 UBL[6] 95 134 VSS n12ll L=6e-08 W=7.5e-07 $X=7835 $Y=30230 $D=0
M150 134 95 UBL[6] VSS n12ll L=6e-08 W=7.5e-07 $X=7835 $Y=30510 $D=0
M151 VSS 136 128 VSS n12ll L=6e-08 W=8e-07 $X=7885 $Y=5385 $D=0
M152 VSS 137 129 VSS n12ll L=6e-08 W=8e-07 $X=7885 $Y=27185 $D=0
M153 VSS 128 133 VSS n12ll L=6e-08 W=1.52e-06 $X=7930 $Y=4590 $D=0
M154 139 145 VSS VSS n12ll L=6e-08 W=1.52e-06 $X=7930 $Y=4860 $D=0
M155 VSS 146 140 VSS n12ll L=6e-08 W=1.52e-06 $X=7930 $Y=28450 $D=0
M156 134 129 VSS VSS n12ll L=6e-08 W=1.52e-06 $X=7930 $Y=28720 $D=0
M157 203 132 VSS VSS n12ll L=6e-08 W=8e-07 $X=8165 $Y=5385 $D=0
M158 204 132 VSS VSS n12ll L=6e-08 W=8e-07 $X=8165 $Y=27185 $D=0
M159 202 126 125 VSS n12ll L=6e-08 W=1e-06 $X=8170 $Y=17700 $D=0
M160 VSS 138 202 VSS n12ll L=6e-08 W=1e-06 $X=8170 $Y=17920 $D=0
M161 135 BWEN VSS VSS n12ll L=6e-08 W=4e-07 $X=8325 $Y=12440 $D=0
M162 136 65 203 VSS n12ll L=6e-08 W=8e-07 $X=8365 $Y=5385 $D=0
M163 137 66 204 VSS n12ll L=6e-08 W=8e-07 $X=8365 $Y=27185 $D=0
M164 138 144 VSS VSS n12ll L=6e-08 W=4e-07 $X=8420 $Y=18820 $D=0
M165 205 SACK1 141 VSS n12ll L=6e-08 W=4e-07 $X=8475 $Y=16120 $D=0
M166 VSS SACK4 205 VSS n12ll L=6e-08 W=4e-07 $X=8695 $Y=16120 $D=0
M167 VSS 144 138 VSS n12ll L=6e-08 W=4e-07 $X=8710 $Y=18820 $D=0
M168 LBL[7] 95 139 VSS n12ll L=6e-08 W=7.5e-07 $X=8775 $Y=2800 $D=0
M169 139 95 LBL[7] VSS n12ll L=6e-08 W=7.5e-07 $X=8775 $Y=3080 $D=0
M170 LBLX[7] 72 139 VSS n12ll L=6e-08 W=7.5e-07 $X=8775 $Y=3360 $D=0
M171 139 72 LBLX[7] VSS n12ll L=6e-08 W=7.5e-07 $X=8775 $Y=3640 $D=0
M172 UBLX[7] 72 140 VSS n12ll L=6e-08 W=7.5e-07 $X=8775 $Y=29670 $D=0
M173 140 72 UBLX[7] VSS n12ll L=6e-08 W=7.5e-07 $X=8775 $Y=29950 $D=0
M174 UBL[7] 95 140 VSS n12ll L=6e-08 W=7.5e-07 $X=8775 $Y=30230 $D=0
M175 140 95 UBL[7] VSS n12ll L=6e-08 W=7.5e-07 $X=8775 $Y=30510 $D=0
M176 206 65 142 VSS n12ll L=6e-08 W=8e-07 $X=8935 $Y=5385 $D=0
M177 207 66 143 VSS n12ll L=6e-08 W=8e-07 $X=8935 $Y=27185 $D=0
M178 VSS VSS BWEN VSS n12ll L=6e-08 W=2e-07 $X=8970 $Y=12475 $D=0
M179 120 141 VSS VSS n12ll L=6e-08 W=5e-07 $X=8985 $Y=16120 $D=0
M180 144 SACK4 VSS VSS n12ll L=6e-08 W=4e-07 $X=9040 $Y=18820 $D=0
M181 VSS 131 206 VSS n12ll L=6e-08 W=8e-07 $X=9135 $Y=5385 $D=0
M182 VSS 131 207 VSS n12ll L=6e-08 W=8e-07 $X=9135 $Y=27185 $D=0
M183 VSS YX[7] 131 VSS n12ll L=6e-08 W=4e-07 $X=9140 $Y=22635 $D=0
M184 132 YX[6] VSS VSS n12ll L=6e-08 W=4e-07 $X=9140 $Y=22925 $D=0
M185 145 142 VSS VSS n12ll L=6e-08 W=8e-07 $X=9415 $Y=5385 $D=0
M186 146 143 VSS VSS n12ll L=6e-08 W=8e-07 $X=9415 $Y=27185 $D=0
M187 59 YX[1] VDD VDD p12ll L=6e-08 W=8e-07 $X=350 $Y=10365 $D=2
M188 LBL[0] 57 VDD VDD p12ll L=6e-08 W=1e-06 $X=375 $Y=1230 $D=2
M189 UBL[0] 58 VDD VDD p12ll L=6e-08 W=1e-06 $X=375 $Y=31140 $D=2
M190 VDD YX[0] 60 VDD p12ll L=6e-08 W=8e-07 $X=400 $Y=22905 $D=2
M191 VDD 63 57 VDD p12ll L=6e-08 W=6e-07 $X=445 $Y=6685 $D=2
M192 VDD 64 58 VDD p12ll L=6e-08 W=6e-07 $X=445 $Y=26085 $D=2
M193 LBLX[0] 57 LBL[0] VDD p12ll L=6e-08 W=1e-06 $X=685 $Y=1230 $D=2
M194 UBLX[0] 58 UBL[0] VDD p12ll L=6e-08 W=1e-06 $X=685 $Y=31140 $D=2
M195 63 60 VDD VDD p12ll L=6e-08 W=6e-07 $X=775 $Y=6685 $D=2
M196 64 60 VDD VDD p12ll L=6e-08 W=6e-07 $X=775 $Y=26085 $D=2
M197 VDD 57 LBLX[0] VDD p12ll L=6e-08 W=1e-06 $X=995 $Y=1230 $D=2
M198 VDD 58 UBLX[0] VDD p12ll L=6e-08 W=1e-06 $X=995 $Y=31140 $D=2
M199 VDD 65 63 VDD p12ll L=6e-08 W=6e-07 $X=1045 $Y=6685 $D=2
M200 VDD 66 64 VDD p12ll L=6e-08 W=6e-07 $X=1045 $Y=26085 $D=2
M201 121 63 LBLX[0] VDD p12ll L=6e-08 W=6e-07 $X=1060 $Y=7885 $D=2
M202 113 63 LBL[0] VDD p12ll L=6e-08 W=6e-07 $X=1060 $Y=8755 $D=2
M203 113 64 UBL[0] VDD p12ll L=6e-08 W=6e-07 $X=1060 $Y=24015 $D=2
M204 121 64 UBLX[0] VDD p12ll L=6e-08 W=6e-07 $X=1060 $Y=24885 $D=2
M205 LBLX[1] 70 121 VDD p12ll L=6e-08 W=6e-07 $X=1360 $Y=7885 $D=2
M206 LBL[1] 70 113 VDD p12ll L=6e-08 W=6e-07 $X=1360 $Y=8755 $D=2
M207 UBL[1] 71 113 VDD p12ll L=6e-08 W=6e-07 $X=1360 $Y=24015 $D=2
M208 UBLX[1] 71 121 VDD p12ll L=6e-08 W=6e-07 $X=1360 $Y=24885 $D=2
M209 70 65 VDD VDD p12ll L=6e-08 W=6e-07 $X=1375 $Y=6685 $D=2
M210 71 66 VDD VDD p12ll L=6e-08 W=6e-07 $X=1375 $Y=26085 $D=2
M211 VDD VDD DATA VDD p12ll L=6e-08 W=2e-07 $X=1410 $Y=15185 $D=2
M212 LBLX[1] 74 VDD VDD p12ll L=6e-08 W=1e-06 $X=1425 $Y=1230 $D=2
M213 UBLX[1] 75 VDD VDD p12ll L=6e-08 W=1e-06 $X=1425 $Y=31140 $D=2
M214 VDD DATA 67 VDD p12ll L=6e-08 W=4e-07 $X=1445 $Y=13450 $D=2
M215 VDD 59 70 VDD p12ll L=6e-08 W=6e-07 $X=1645 $Y=6685 $D=2
M216 VDD 59 71 VDD p12ll L=6e-08 W=6e-07 $X=1645 $Y=26085 $D=2
M217 LBL[1] 74 LBLX[1] VDD p12ll L=6e-08 W=1e-06 $X=1735 $Y=1230 $D=2
M218 UBL[1] 75 UBLX[1] VDD p12ll L=6e-08 W=1e-06 $X=1735 $Y=31140 $D=2
M219 72 77 VDD VDD p12ll L=6e-08 W=2e-06 $X=1790 $Y=19770 $D=2
M220 76 67 VDD VDD p12ll L=3e-07 W=4e-07 $X=1835 $Y=13450 $D=2
M221 73 91 VDD VDD p12ll L=6e-08 W=4e-07 $X=1860 $Y=14985 $D=2
M222 74 70 VDD VDD p12ll L=6e-08 W=6e-07 $X=1975 $Y=6685 $D=2
M223 75 71 VDD VDD p12ll L=6e-08 W=6e-07 $X=1975 $Y=26085 $D=2
M224 VDD 74 LBL[1] VDD p12ll L=6e-08 W=1e-06 $X=2045 $Y=1230 $D=2
M225 VDD 75 UBL[1] VDD p12ll L=6e-08 W=1e-06 $X=2045 $Y=31140 $D=2
M226 VDD 77 72 VDD p12ll L=6e-08 W=2e-06 $X=2080 $Y=19770 $D=2
M227 77 73 VDD VDD p12ll L=6e-08 W=8e-07 $X=2415 $Y=19770 $D=2
M228 VDD 83 80 VDD p12ll L=6e-08 W=1e-06 $X=2510 $Y=14420 $D=2
M229 VDD 80 77 VDD p12ll L=6e-08 W=8e-07 $X=2705 $Y=19770 $D=2
M230 83 WE VDD VDD p12ll L=6e-08 W=4e-07 $X=2800 $Y=15020 $D=2
M231 VDD 76 84 VDD p12ll L=2e-07 W=4e-07 $X=2845 $Y=13460 $D=2
M232 LBL[2] 78 VDD VDD p12ll L=6e-08 W=1e-06 $X=2855 $Y=1230 $D=2
M233 UBL[2] 79 VDD VDD p12ll L=6e-08 W=1e-06 $X=2855 $Y=31140 $D=2
M234 VDD 87 78 VDD p12ll L=6e-08 W=6e-07 $X=2925 $Y=6685 $D=2
M235 VDD 88 79 VDD p12ll L=6e-08 W=6e-07 $X=2925 $Y=26085 $D=2
M236 VDD 101 83 VDD p12ll L=6e-08 W=4e-07 $X=3090 $Y=15020 $D=2
M237 LBLX[2] 78 LBL[2] VDD p12ll L=6e-08 W=1e-06 $X=3165 $Y=1230 $D=2
M238 UBLX[2] 79 UBL[2] VDD p12ll L=6e-08 W=1e-06 $X=3165 $Y=31140 $D=2
M239 90 80 VDD VDD p12ll L=6e-08 W=8e-07 $X=3185 $Y=19770 $D=2
M240 87 82 VDD VDD p12ll L=6e-08 W=6e-07 $X=3255 $Y=6685 $D=2
M241 88 82 VDD VDD p12ll L=6e-08 W=6e-07 $X=3255 $Y=26085 $D=2
M242 89 84 VDD VDD p12ll L=6e-08 W=7e-07 $X=3355 $Y=13385 $D=2
M243 VDD 91 94 VDD p12ll L=3e-07 W=1.2e-07 $X=3460 $Y=14605 $D=2
M244 VDD 78 LBLX[2] VDD p12ll L=6e-08 W=1e-06 $X=3475 $Y=1230 $D=2
M245 VDD 91 90 VDD p12ll L=6e-08 W=8e-07 $X=3475 $Y=19770 $D=2
M246 VDD 79 UBLX[2] VDD p12ll L=6e-08 W=1e-06 $X=3475 $Y=31140 $D=2
M247 VDD 65 87 VDD p12ll L=6e-08 W=6e-07 $X=3525 $Y=6685 $D=2
M248 VDD 66 88 VDD p12ll L=6e-08 W=6e-07 $X=3525 $Y=26085 $D=2
M249 121 87 LBLX[2] VDD p12ll L=6e-08 W=6e-07 $X=3540 $Y=7885 $D=2
M250 113 87 LBL[2] VDD p12ll L=6e-08 W=6e-07 $X=3540 $Y=8755 $D=2
M251 113 88 UBL[2] VDD p12ll L=6e-08 W=6e-07 $X=3540 $Y=24015 $D=2
M252 121 88 UBLX[2] VDD p12ll L=6e-08 W=6e-07 $X=3540 $Y=24885 $D=2
M253 94 CLK 89 VDD p12ll L=6e-08 W=7e-07 $X=3700 $Y=13385 $D=2
M254 95 90 VDD VDD p12ll L=6e-08 W=2e-06 $X=3805 $Y=19770 $D=2
M255 VDD YX[2] 82 VDD p12ll L=6e-08 W=8e-07 $X=3810 $Y=10455 $D=2
M256 81 YX[3] VDD VDD p12ll L=6e-08 W=8e-07 $X=3810 $Y=10745 $D=2
M257 LBLX[3] 96 121 VDD p12ll L=6e-08 W=6e-07 $X=3840 $Y=7885 $D=2
M258 LBL[3] 96 113 VDD p12ll L=6e-08 W=6e-07 $X=3840 $Y=8755 $D=2
M259 UBL[3] 97 113 VDD p12ll L=6e-08 W=6e-07 $X=3840 $Y=24015 $D=2
M260 UBLX[3] 97 121 VDD p12ll L=6e-08 W=6e-07 $X=3840 $Y=24885 $D=2
M261 96 65 VDD VDD p12ll L=6e-08 W=6e-07 $X=3855 $Y=6685 $D=2
M262 97 66 VDD VDD p12ll L=6e-08 W=6e-07 $X=3855 $Y=26085 $D=2
M263 LBLX[3] 98 VDD VDD p12ll L=6e-08 W=1e-06 $X=3905 $Y=1230 $D=2
M264 UBLX[3] 99 VDD VDD p12ll L=6e-08 W=1e-06 $X=3905 $Y=31140 $D=2
M265 VDD 90 95 VDD p12ll L=6e-08 W=2e-06 $X=4095 $Y=19770 $D=2
M266 VDD 81 96 VDD p12ll L=6e-08 W=6e-07 $X=4125 $Y=6685 $D=2
M267 VDD 81 97 VDD p12ll L=6e-08 W=6e-07 $X=4125 $Y=26085 $D=2
M268 LBL[3] 98 LBLX[3] VDD p12ll L=6e-08 W=1e-06 $X=4215 $Y=1230 $D=2
M269 UBL[3] 99 UBLX[3] VDD p12ll L=6e-08 W=1e-06 $X=4215 $Y=31140 $D=2
M270 98 96 VDD VDD p12ll L=6e-08 W=6e-07 $X=4455 $Y=6685 $D=2
M271 99 97 VDD VDD p12ll L=6e-08 W=6e-07 $X=4455 $Y=26085 $D=2
M272 VDD 94 91 VDD p12ll L=6e-08 W=8e-07 $X=4485 $Y=13370 $D=2
M273 VDD 98 LBL[3] VDD p12ll L=6e-08 W=1e-06 $X=4525 $Y=1230 $D=2
M274 VDD 99 UBL[3] VDD p12ll L=6e-08 W=1e-06 $X=4525 $Y=31140 $D=2
M275 VDD 109 DOUT VDD p12ll L=6e-08 W=1e-06 $X=4675 $Y=14425 $D=2
M276 110 101 VDD VDD p12ll L=3e-07 W=1.2e-07 $X=4865 $Y=13890 $D=2
M277 DOUT 109 VDD VDD p12ll L=6e-08 W=1e-06 $X=4965 $Y=14425 $D=2
M278 113 120 100 VDD p12ll L=6e-08 W=1.4e-06 $X=5080 $Y=20430 $D=2
M279 VDD 109 DOUT VDD p12ll L=6e-08 W=1e-06 $X=5255 $Y=14425 $D=2
M280 VDD YX[4] 105 VDD p12ll L=6e-08 W=8e-07 $X=5315 $Y=10330 $D=2
M281 65 AS VDD VDD p12ll L=6e-08 W=8e-07 $X=5315 $Y=10630 $D=2
M282 LBL[4] 103 VDD VDD p12ll L=6e-08 W=1e-06 $X=5335 $Y=1230 $D=2
M283 UBL[4] 104 VDD VDD p12ll L=6e-08 W=1e-06 $X=5335 $Y=31140 $D=2
M284 VDD 110 101 VDD p12ll L=6e-08 W=4e-07 $X=5345 $Y=13290 $D=2
M285 VDD 111 103 VDD p12ll L=6e-08 W=6e-07 $X=5405 $Y=6685 $D=2
M286 VDD 112 104 VDD p12ll L=6e-08 W=6e-07 $X=5405 $Y=26085 $D=2
M287 108 100 VDD VDD p12ll L=1e-07 W=4e-07 $X=5460 $Y=19765 $D=2
M288 109 100 VDD VDD p12ll L=6e-08 W=1e-06 $X=5545 $Y=14425 $D=2
M289 LBLX[4] 103 LBL[4] VDD p12ll L=6e-08 W=1e-06 $X=5645 $Y=1230 $D=2
M290 UBLX[4] 104 UBL[4] VDD p12ll L=6e-08 W=1e-06 $X=5645 $Y=31140 $D=2
M291 111 105 VDD VDD p12ll L=6e-08 W=6e-07 $X=5735 $Y=6685 $D=2
M292 112 105 VDD VDD p12ll L=6e-08 W=6e-07 $X=5735 $Y=26085 $D=2
M293 VDD 119 109 VDD p12ll L=6e-08 W=1e-06 $X=5835 $Y=14425 $D=2
M294 113 138 VDD VDD p12ll L=6e-08 W=1e-06 $X=5880 $Y=20750 $D=2
M295 VDD 100 108 VDD p12ll L=1e-07 W=4e-07 $X=5920 $Y=19765 $D=2
M296 VDD 103 LBLX[4] VDD p12ll L=6e-08 W=1e-06 $X=5955 $Y=1230 $D=2
M297 VDD 104 UBLX[4] VDD p12ll L=6e-08 W=1e-06 $X=5955 $Y=31140 $D=2
M298 VDD 65 111 VDD p12ll L=6e-08 W=6e-07 $X=6005 $Y=6685 $D=2
M299 VDD 66 112 VDD p12ll L=6e-08 W=6e-07 $X=6005 $Y=26085 $D=2
M300 121 111 LBLX[4] VDD p12ll L=6e-08 W=6e-07 $X=6020 $Y=7885 $D=2
M301 113 111 LBL[4] VDD p12ll L=6e-08 W=6e-07 $X=6020 $Y=8755 $D=2
M302 113 112 UBL[4] VDD p12ll L=6e-08 W=6e-07 $X=6020 $Y=24015 $D=2
M303 121 112 UBLX[4] VDD p12ll L=6e-08 W=6e-07 $X=6020 $Y=24885 $D=2
M304 114 CLK 110 VDD p12ll L=6e-08 W=7e-07 $X=6120 $Y=13300 $D=2
M305 121 138 113 VDD p12ll L=6e-08 W=1e-06 $X=6170 $Y=20750 $D=2
M306 VDD AXS 66 VDD p12ll L=6e-08 W=8e-07 $X=6265 $Y=22645 $D=2
M307 102 YX[5] VDD VDD p12ll L=6e-08 W=8e-07 $X=6265 $Y=22990 $D=2
M308 LBLX[5] 117 121 VDD p12ll L=6e-08 W=6e-07 $X=6320 $Y=7885 $D=2
M309 LBL[5] 117 113 VDD p12ll L=6e-08 W=6e-07 $X=6320 $Y=8755 $D=2
M310 UBL[5] 118 113 VDD p12ll L=6e-08 W=6e-07 $X=6320 $Y=24015 $D=2
M311 UBLX[5] 118 121 VDD p12ll L=6e-08 W=6e-07 $X=6320 $Y=24885 $D=2
M312 117 65 VDD VDD p12ll L=6e-08 W=6e-07 $X=6335 $Y=6685 $D=2
M313 118 66 VDD VDD p12ll L=6e-08 W=6e-07 $X=6335 $Y=26085 $D=2
M314 100 108 VDD VDD p12ll L=1e-07 W=4e-07 $X=6380 $Y=19765 $D=2
M315 LBLX[5] 123 VDD VDD p12ll L=6e-08 W=1e-06 $X=6385 $Y=1230 $D=2
M316 UBLX[5] 124 VDD VDD p12ll L=6e-08 W=1e-06 $X=6385 $Y=31140 $D=2
M317 VDD 138 121 VDD p12ll L=6e-08 W=1e-06 $X=6460 $Y=20750 $D=2
M318 VDD 122 114 VDD p12ll L=6e-08 W=7e-07 $X=6490 $Y=13300 $D=2
M319 119 109 VDD VDD p12ll L=6e-08 W=1e-06 $X=6515 $Y=14425 $D=2
M320 VDD 102 117 VDD p12ll L=6e-08 W=6e-07 $X=6605 $Y=6685 $D=2
M321 VDD 102 118 VDD p12ll L=6e-08 W=6e-07 $X=6605 $Y=26085 $D=2
M322 LBL[5] 123 LBLX[5] VDD p12ll L=6e-08 W=1e-06 $X=6695 $Y=1230 $D=2
M323 UBL[5] 124 UBLX[5] VDD p12ll L=6e-08 W=1e-06 $X=6695 $Y=31140 $D=2
M324 VDD 108 119 VDD p12ll L=6e-08 W=1e-06 $X=6805 $Y=14425 $D=2
M325 122 127 VDD VDD p12ll L=2e-07 W=4e-07 $X=6830 $Y=13565 $D=2
M326 VDD 108 100 VDD p12ll L=1e-07 W=4e-07 $X=6840 $Y=19765 $D=2
M327 123 117 VDD VDD p12ll L=6e-08 W=6e-07 $X=6935 $Y=6685 $D=2
M328 124 118 VDD VDD p12ll L=6e-08 W=6e-07 $X=6935 $Y=26085 $D=2
M329 VDD 123 LBL[5] VDD p12ll L=6e-08 W=1e-06 $X=7005 $Y=1230 $D=2
M330 VDD 124 UBL[5] VDD p12ll L=6e-08 W=1e-06 $X=7005 $Y=31140 $D=2
M331 108 120 121 VDD p12ll L=6e-08 W=1.4e-06 $X=7260 $Y=20430 $D=2
M332 VDD 130 126 VDD p12ll L=6e-08 W=1e-06 $X=7465 $Y=14395 $D=2
M333 VDD 135 127 VDD p12ll L=3e-07 W=4e-07 $X=7735 $Y=13450 $D=2
M334 130 SACK1 VDD VDD p12ll L=6e-08 W=4e-07 $X=7755 $Y=14995 $D=2
M335 LBL[6] 128 VDD VDD p12ll L=6e-08 W=1e-06 $X=7815 $Y=1230 $D=2
M336 UBL[6] 129 VDD VDD p12ll L=6e-08 W=1e-06 $X=7815 $Y=31140 $D=2
M337 VDD YX[7] 131 VDD p12ll L=6e-08 W=8e-07 $X=7850 $Y=22635 $D=2
M338 132 YX[6] VDD VDD p12ll L=6e-08 W=8e-07 $X=7850 $Y=22925 $D=2
M339 VDD 136 128 VDD p12ll L=6e-08 W=6e-07 $X=7885 $Y=6685 $D=2
M340 VDD 137 129 VDD p12ll L=6e-08 W=6e-07 $X=7885 $Y=26085 $D=2
M341 LBLX[6] 128 LBL[6] VDD p12ll L=6e-08 W=1e-06 $X=8125 $Y=1230 $D=2
M342 UBLX[6] 129 UBL[6] VDD p12ll L=6e-08 W=1e-06 $X=8125 $Y=31140 $D=2
M343 136 132 VDD VDD p12ll L=6e-08 W=6e-07 $X=8215 $Y=6685 $D=2
M344 137 132 VDD VDD p12ll L=6e-08 W=6e-07 $X=8215 $Y=26085 $D=2
M345 135 BWEN VDD VDD p12ll L=6e-08 W=4e-07 $X=8325 $Y=13450 $D=2
M346 141 SACK1 VDD VDD p12ll L=6e-08 W=4e-07 $X=8405 $Y=14990 $D=2
M347 138 144 VDD VDD p12ll L=6e-08 W=8e-07 $X=8420 $Y=19840 $D=2
M348 VDD 128 LBLX[6] VDD p12ll L=6e-08 W=1e-06 $X=8435 $Y=1230 $D=2
M349 VDD 129 UBLX[6] VDD p12ll L=6e-08 W=1e-06 $X=8435 $Y=31140 $D=2
M350 VDD 65 136 VDD p12ll L=6e-08 W=6e-07 $X=8485 $Y=6685 $D=2
M351 VDD 66 137 VDD p12ll L=6e-08 W=6e-07 $X=8485 $Y=26085 $D=2
M352 121 136 LBLX[6] VDD p12ll L=6e-08 W=6e-07 $X=8500 $Y=7885 $D=2
M353 113 136 LBL[6] VDD p12ll L=6e-08 W=6e-07 $X=8500 $Y=8755 $D=2
M354 113 137 UBL[6] VDD p12ll L=6e-08 W=6e-07 $X=8500 $Y=24015 $D=2
M355 121 137 UBLX[6] VDD p12ll L=6e-08 W=6e-07 $X=8500 $Y=24885 $D=2
M356 VDD SACK4 141 VDD p12ll L=6e-08 W=4e-07 $X=8695 $Y=14990 $D=2
M357 VDD 144 138 VDD p12ll L=6e-08 W=8e-07 $X=8710 $Y=19840 $D=2
M358 LBLX[7] 142 121 VDD p12ll L=6e-08 W=6e-07 $X=8800 $Y=7885 $D=2
M359 LBL[7] 142 113 VDD p12ll L=6e-08 W=6e-07 $X=8800 $Y=8755 $D=2
M360 UBL[7] 143 113 VDD p12ll L=6e-08 W=6e-07 $X=8800 $Y=24015 $D=2
M361 UBLX[7] 143 121 VDD p12ll L=6e-08 W=6e-07 $X=8800 $Y=24885 $D=2
M362 142 65 VDD VDD p12ll L=6e-08 W=6e-07 $X=8815 $Y=6685 $D=2
M363 143 66 VDD VDD p12ll L=6e-08 W=6e-07 $X=8815 $Y=26085 $D=2
M364 LBLX[7] 145 VDD VDD p12ll L=6e-08 W=1e-06 $X=8865 $Y=1230 $D=2
M365 UBLX[7] 146 VDD VDD p12ll L=6e-08 W=1e-06 $X=8865 $Y=31140 $D=2
M366 VDD VDD BWEN VDD p12ll L=6e-08 W=2e-07 $X=8970 $Y=13520 $D=2
M367 120 141 VDD VDD p12ll L=6e-08 W=1e-06 $X=8985 $Y=14390 $D=2
M368 144 SACK4 VDD VDD p12ll L=6e-08 W=8e-07 $X=9040 $Y=19840 $D=2
M369 VDD 131 142 VDD p12ll L=6e-08 W=6e-07 $X=9085 $Y=6685 $D=2
M370 VDD 131 143 VDD p12ll L=6e-08 W=6e-07 $X=9085 $Y=26085 $D=2
M371 LBL[7] 145 LBLX[7] VDD p12ll L=6e-08 W=1e-06 $X=9175 $Y=1230 $D=2
M372 UBL[7] 146 UBLX[7] VDD p12ll L=6e-08 W=1e-06 $X=9175 $Y=31140 $D=2
M373 145 142 VDD VDD p12ll L=6e-08 W=6e-07 $X=9415 $Y=6685 $D=2
M374 146 143 VDD VDD p12ll L=6e-08 W=6e-07 $X=9415 $Y=26085 $D=2
M375 VDD 145 LBL[7] VDD p12ll L=6e-08 W=1e-06 $X=9485 $Y=1230 $D=2
M376 VDD 146 UBL[7] VDD p12ll L=6e-08 W=1e-06 $X=9485 $Y=31140 $D=2
.ENDS
***************************************
.SUBCKT Y8_X128_D1_BW_620_VHSSP 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149
** N=186 EP=149 IP=225 FDC=6905
X0 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170
+ Y8_X64_1_DOWN_BW_620_VHSSP $T=0 41705 1 0 $X=-1320 $Y=0
X1 1 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108
+ 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128
+ 129 130 131 132 133 134 2 171 172 173 174 175 176 177 178 179 180 181 182 183
+ 184 185 186
+ Y8_X64_1_UP_620_VHSSP $T=0 75080 0 0 $X=-1320 $Y=74385
X2 1 2 155 171 156 172 140 149 67 157 173 158 174 142 159 175 137 160 176 138
+ 136 161 177 162 178 141 148 68 163 179 145 164 180 144 165 181 166 182 167 183
+ 147 168 184 139 143 169 185 170 186 135 69 146
+ YMX8SAWR_BW_620 $T=0 41705 0 0 $X=-520 $Y=41330
.ENDS
***************************************
.SUBCKT Y8_X128_D2_BW_620_VHSSP 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152
** N=158 EP=152 IP=308 FDC=13810
X0 1 2 66 65 64 63 62 61 60 59 58 57 56 55 54 53 52 51 50 49
+ 48 47 46 45 44 43 42 41 40 39 38 37 36 35 34 33 32 31 30 29
+ 28 27 26 25 24 23 22 21 20 19 18 17 16 15 14 13 12 11 10 9
+ 8 7 6 5 4 3 132 133 134 67 68 69 70 71 72 73 74 75 76 77
+ 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97
+ 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117
+ 118 119 120 121 122 123 124 125 126 127 128 129 130 131 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152
+ Y8_X128_D1_BW_620_VHSSP $T=0 0 0 0 $X=-1320 $Y=0
X1 1 2 66 65 64 63 62 61 60 59 58 57 56 55 54 53 52 51 50 49
+ 48 47 46 45 44 43 42 41 40 39 38 37 36 35 34 33 32 31 30 29
+ 28 27 26 25 24 23 22 21 20 19 18 17 16 15 14 13 12 11 10 9
+ 8 7 6 5 4 3 135 136 137 67 68 69 70 71 72 73 74 75 76 77
+ 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97
+ 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117
+ 118 119 120 121 122 123 124 125 126 127 128 129 130 131 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152
+ Y8_X128_D1_BW_620_VHSSP $T=19840 0 1 180 $X=8600 $Y=0
.ENDS
***************************************
.SUBCKT 65smic_062swl_svt_dummycell_v0p0_st 1 2 3 4 5
** N=10 EP=5 IP=0 FDC=6
M0 3 1 7 2 DNNPGSVT L=7.5e-08 W=1.25e-07 $X=150 $Y=335 $D=96
M1 8 2 5 2 DNNPGSVT L=7.5e-08 W=1.25e-07 $X=965 $Y=90 $D=96
M2 7 8 2 2 DNNPDSVT L=6.5e-08 W=2.1e-07 $X=125 $Y=90 $D=95
M3 2 7 8 2 DNNPDSVT L=6.5e-08 W=2.1e-07 $X=905 $Y=345 $D=95
M4 7 8 4 4 DNPLSVT L=6.5e-08 W=9.5e-08 $X=470 $Y=90 $D=97
M5 4 7 8 4 DNPLSVT L=6.5e-08 W=9.5e-08 $X=675 $Y=345 $D=97
.ENDS
***************************************
.SUBCKT bitcell_dummy_left_2A_st_620_VHSSP 1 2 3 4 5
** N=7 EP=5 IP=12 FDC=12
X0 1 2 7 3 4 65smic_062swl_svt_dummycell_v0p0_st $T=0 0 0 0 $X=-125 $Y=-185
X1 5 2 7 3 4 65smic_062swl_svt_dummycell_v0p0_st $T=0 1000 1 0 $X=-125 $Y=315
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4 5 6 7
** N=8 EP=7 IP=12 FDC=24
X0 1 3 4 5 2 bitcell_dummy_left_2A_st_620_VHSSP $T=0 -1000 0 0 $X=-125 $Y=-1185
X1 6 3 4 5 7 bitcell_dummy_left_2A_st_620_VHSSP $T=0 0 0 0 $X=-125 $Y=-185
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8 9 10 11
** N=12 EP=11 IP=16 FDC=48
X0 2 3 1 6 7 4 5 ICV_7 $T=0 -2000 0 0 $X=-125 $Y=-3185
X1 8 9 1 6 7 10 11 ICV_7 $T=0 0 0 0 $X=-125 $Y=-1185
.ENDS
***************************************
.SUBCKT bitcell_dummy_left_2B_st_620_VHSSP 1 2 3 4 5 6 7
** N=8 EP=7 IP=12 FDC=12
X0 1 2 3 4 5 65smic_062swl_svt_dummycell_v0p0_st $T=0 500 1 0 $X=-125 $Y=-185
X1 6 2 7 4 5 65smic_062swl_svt_dummycell_v0p0_st $T=0 500 0 0 $X=-125 $Y=315
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6 7 8 10
** N=11 EP=9 IP=16 FDC=24
X0 2 1 4 5 10 3 11 bitcell_dummy_left_2B_st_620_VHSSP $T=0 -1000 0 0 $X=-125 $Y=-1185
X1 6 1 11 5 10 7 8 bitcell_dummy_left_2B_st_620_VHSSP $T=0 0 0 0 $X=-125 $Y=-185
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5 6 7 8 9 10 11 12 14
** N=15 EP=13 IP=20 FDC=48
X0 1 2 3 6 7 4 5 15 14 ICV_9 $T=0 -2000 0 0 $X=-125 $Y=-3185
X1 1 8 9 15 7 10 11 12 14 ICV_9 $T=0 0 0 0 $X=-125 $Y=-1185
.ENDS
***************************************
.SUBCKT LEAF_XDEC_TOP_POWER_VHS
** N=37 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VDD VSS
.ENDS
***************************************
.SUBCKT LEAF_XDEC4_VHSSRAM VDD 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 VSS 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78
** N=228 EP=78 IP=0 FDC=792
M0 2 105 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=695 $D=0
M1 VSS 105 2 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=945 $D=0
M2 3 106 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=1195 $D=0
M3 VSS 106 3 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=1445 $D=0
M4 4 107 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=1695 $D=0
M5 VSS 107 4 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=1945 $D=0
M6 5 108 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=2195 $D=0
M7 VSS 108 5 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=2445 $D=0
M8 6 109 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=2695 $D=0
M9 VSS 109 6 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=2945 $D=0
M10 7 110 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=3195 $D=0
M11 VSS 110 7 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=3445 $D=0
M12 8 111 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=3695 $D=0
M13 VSS 111 8 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=3945 $D=0
M14 9 112 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=4195 $D=0
M15 VSS 112 9 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=4445 $D=0
M16 10 113 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=4695 $D=0
M17 VSS 113 10 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=4945 $D=0
M18 11 114 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=5195 $D=0
M19 VSS 114 11 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=5445 $D=0
M20 12 115 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=5695 $D=0
M21 VSS 115 12 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=5945 $D=0
M22 13 116 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=6195 $D=0
M23 VSS 116 13 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=6445 $D=0
M24 14 117 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=6695 $D=0
M25 VSS 117 14 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=6945 $D=0
M26 15 118 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=7195 $D=0
M27 VSS 118 15 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=7445 $D=0
M28 16 119 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=7695 $D=0
M29 VSS 119 16 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=7945 $D=0
M30 17 120 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=8195 $D=0
M31 VSS 120 17 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=8445 $D=0
M32 18 121 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=8695 $D=0
M33 VSS 121 18 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=8945 $D=0
M34 19 122 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=9195 $D=0
M35 VSS 122 19 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=9445 $D=0
M36 20 123 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=9695 $D=0
M37 VSS 123 20 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=9945 $D=0
M38 21 124 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=10195 $D=0
M39 VSS 124 21 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=10445 $D=0
M40 22 125 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=10695 $D=0
M41 VSS 125 22 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=10945 $D=0
M42 23 126 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=11195 $D=0
M43 VSS 126 23 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=11445 $D=0
M44 24 127 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=11695 $D=0
M45 VSS 127 24 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=11945 $D=0
M46 25 128 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=12195 $D=0
M47 VSS 128 25 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=12445 $D=0
M48 26 129 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=12695 $D=0
M49 VSS 129 26 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=12945 $D=0
M50 27 130 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=13195 $D=0
M51 VSS 130 27 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=13445 $D=0
M52 28 131 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=13695 $D=0
M53 VSS 131 28 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=13945 $D=0
M54 29 132 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=14195 $D=0
M55 VSS 132 29 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=14445 $D=0
M56 30 133 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=14695 $D=0
M57 VSS 133 30 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=14945 $D=0
M58 31 134 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=15195 $D=0
M59 VSS 134 31 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=15445 $D=0
M60 32 135 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=15695 $D=0
M61 VSS 135 32 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=15945 $D=0
M62 33 136 VSS VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=16195 $D=0
M63 VSS 136 33 VSS n12ll L=6e-08 W=1e-06 $X=3890 $Y=16445 $D=0
M64 105 137 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=695 $D=0
M65 VSS 137 105 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=945 $D=0
M66 105 137 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=1195 $D=0
M67 VSS 137 105 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=1445 $D=0
M68 106 138 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=1695 $D=0
M69 VSS 138 106 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=1945 $D=0
M70 106 138 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=2195 $D=0
M71 VSS 138 106 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=2445 $D=0
M72 107 139 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=2695 $D=0
M73 VSS 139 107 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=2945 $D=0
M74 107 139 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=3195 $D=0
M75 VSS 139 107 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=3445 $D=0
M76 108 140 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=3695 $D=0
M77 VSS 140 108 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=3945 $D=0
M78 108 140 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=4195 $D=0
M79 VSS 140 108 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=4445 $D=0
M80 117 141 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=4695 $D=0
M81 VSS 141 117 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=4945 $D=0
M82 117 141 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=5195 $D=0
M83 VSS 141 117 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=5445 $D=0
M84 118 142 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=5695 $D=0
M85 VSS 142 118 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=5945 $D=0
M86 118 142 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=6195 $D=0
M87 VSS 142 118 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=6445 $D=0
M88 119 143 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=6695 $D=0
M89 VSS 143 119 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=6945 $D=0
M90 119 143 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=7195 $D=0
M91 VSS 143 119 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=7445 $D=0
M92 120 144 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=7695 $D=0
M93 VSS 144 120 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=7945 $D=0
M94 120 144 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=8195 $D=0
M95 VSS 144 120 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=8445 $D=0
M96 121 145 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=8695 $D=0
M97 VSS 145 121 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=8945 $D=0
M98 121 145 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=9195 $D=0
M99 VSS 145 121 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=9445 $D=0
M100 122 146 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=9695 $D=0
M101 VSS 146 122 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=9945 $D=0
M102 122 146 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=10195 $D=0
M103 VSS 146 122 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=10445 $D=0
M104 123 147 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=10695 $D=0
M105 VSS 147 123 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=10945 $D=0
M106 123 147 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=11195 $D=0
M107 VSS 147 123 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=11445 $D=0
M108 124 148 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=11695 $D=0
M109 VSS 148 124 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=11945 $D=0
M110 124 148 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=12195 $D=0
M111 VSS 148 124 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=12445 $D=0
M112 133 149 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=12695 $D=0
M113 VSS 149 133 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=12945 $D=0
M114 133 149 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=13195 $D=0
M115 VSS 149 133 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=13445 $D=0
M116 134 150 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=13695 $D=0
M117 VSS 150 134 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=13945 $D=0
M118 134 150 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=14195 $D=0
M119 VSS 150 134 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=14445 $D=0
M120 135 151 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=14695 $D=0
M121 VSS 151 135 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=14945 $D=0
M122 135 151 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=15195 $D=0
M123 VSS 151 135 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=15445 $D=0
M124 136 152 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=15695 $D=0
M125 VSS 152 136 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=15945 $D=0
M126 136 152 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=16195 $D=0
M127 VSS 152 136 VSS n12ll L=6e-08 W=7.5e-07 $X=5800 $Y=16445 $D=0
M128 137 153 VSS VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=700 $D=0
M129 VSS 154 138 VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=2440 $D=0
M130 139 155 VSS VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=2700 $D=0
M131 VSS 156 140 VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=4440 $D=0
M132 141 157 VSS VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=4700 $D=0
M133 VSS 158 142 VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=6440 $D=0
M134 143 159 VSS VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=6700 $D=0
M135 VSS 160 144 VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=8440 $D=0
M136 145 161 VSS VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=8700 $D=0
M137 VSS 162 146 VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=10440 $D=0
M138 147 163 VSS VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=10700 $D=0
M139 VSS 164 148 VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=12440 $D=0
M140 149 165 VSS VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=12700 $D=0
M141 VSS 166 150 VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=14440 $D=0
M142 151 167 VSS VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=14700 $D=0
M143 VSS 168 152 VSS n12ll L=6e-08 W=8e-07 $X=9870 $Y=16440 $D=0
M144 153 173 35 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=1285 $D=0
M145 36 173 154 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=1855 $D=0
M146 155 173 37 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=3285 $D=0
M147 38 173 156 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=3855 $D=0
M148 157 174 38 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=5285 $D=0
M149 37 174 158 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=5855 $D=0
M150 159 174 36 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=7285 $D=0
M151 35 174 160 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=7855 $D=0
M152 161 175 35 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=9285 $D=0
M153 36 175 162 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=9855 $D=0
M154 163 175 37 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=11285 $D=0
M155 38 175 164 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=11855 $D=0
M156 165 176 38 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=13285 $D=0
M157 37 176 166 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=13855 $D=0
M158 167 176 36 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=15285 $D=0
M159 35 176 168 VSS n12ll L=6e-08 W=6e-07 $X=10020 $Y=15855 $D=0
M160 221 39 VSS VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=3430 $D=0
M161 222 40 221 VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=3720 $D=0
M162 169 VDD 222 VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=4010 $D=0
M163 223 VDD 170 VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=5130 $D=0
M164 224 40 223 VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=5420 $D=0
M165 VSS 41 224 VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=5710 $D=0
M166 225 39 VSS VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=11430 $D=0
M167 226 42 225 VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=11720 $D=0
M168 171 VDD 226 VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=12010 $D=0
M169 227 VDD 172 VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=13130 $D=0
M170 228 42 227 VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=13420 $D=0
M171 VSS 41 228 VSS n12ll L=6e-08 W=8e-07 $X=12695 $Y=13710 $D=0
M172 177 173 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=1120 $D=0
M173 VSS 173 177 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=1405 $D=0
M174 177 173 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=1695 $D=0
M175 VSS 173 177 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=1985 $D=0
M176 173 169 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=2275 $D=0
M177 VSS 169 173 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=2560 $D=0
M178 173 169 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=2850 $D=0
M179 VSS 169 173 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=3140 $D=0
M180 174 170 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=6000 $D=0
M181 VSS 170 174 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=6290 $D=0
M182 174 170 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=6580 $D=0
M183 VSS 170 174 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=6865 $D=0
M184 178 174 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=7155 $D=0
M185 VSS 174 178 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=7445 $D=0
M186 178 174 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=7735 $D=0
M187 VSS 174 178 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=8020 $D=0
M188 179 175 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=9120 $D=0
M189 VSS 175 179 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=9405 $D=0
M190 179 175 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=9695 $D=0
M191 VSS 175 179 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=9985 $D=0
M192 175 171 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=10275 $D=0
M193 VSS 171 175 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=10560 $D=0
M194 175 171 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=10850 $D=0
M195 VSS 171 175 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=11140 $D=0
M196 176 172 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=14000 $D=0
M197 VSS 172 176 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=14290 $D=0
M198 176 172 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=14580 $D=0
M199 VSS 172 176 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=14865 $D=0
M200 180 176 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=15155 $D=0
M201 VSS 176 180 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=15445 $D=0
M202 180 176 VSS VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=15735 $D=0
M203 VSS 176 180 VSS n12ll L=6e-08 W=5e-07 $X=12815 $Y=16020 $D=0
M204 197 181 VSS VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=700 $D=0
M205 VSS 182 198 VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=2440 $D=0
M206 199 183 VSS VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=2700 $D=0
M207 VSS 184 200 VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=4440 $D=0
M208 201 185 VSS VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=4700 $D=0
M209 VSS 186 202 VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=6440 $D=0
M210 203 187 VSS VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=6700 $D=0
M211 VSS 188 204 VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=8440 $D=0
M212 205 189 VSS VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=8700 $D=0
M213 VSS 190 206 VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=10440 $D=0
M214 207 191 VSS VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=10700 $D=0
M215 VSS 192 208 VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=12440 $D=0
M216 209 193 VSS VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=12700 $D=0
M217 VSS 194 210 VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=14440 $D=0
M218 211 195 VSS VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=14700 $D=0
M219 VSS 196 212 VSS n12ll L=6e-08 W=8e-07 $X=16550 $Y=16440 $D=0
M220 181 173 43 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=1290 $D=0
M221 44 173 182 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=1850 $D=0
M222 183 173 45 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=3290 $D=0
M223 46 173 184 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=3850 $D=0
M224 185 174 46 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=5290 $D=0
M225 45 174 186 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=5850 $D=0
M226 187 174 44 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=7290 $D=0
M227 43 174 188 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=7850 $D=0
M228 189 175 43 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=9290 $D=0
M229 44 175 190 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=9850 $D=0
M230 191 175 45 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=11290 $D=0
M231 46 175 192 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=11850 $D=0
M232 193 176 46 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=13290 $D=0
M233 45 176 194 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=13850 $D=0
M234 195 176 44 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=15290 $D=0
M235 43 176 196 VSS n12ll L=6e-08 W=6e-07 $X=16630 $Y=15850 $D=0
M236 109 197 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=695 $D=0
M237 VSS 197 109 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=945 $D=0
M238 109 197 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=1195 $D=0
M239 VSS 197 109 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=1445 $D=0
M240 110 198 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=1695 $D=0
M241 VSS 198 110 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=1945 $D=0
M242 110 198 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=2195 $D=0
M243 VSS 198 110 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=2445 $D=0
M244 111 199 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=2695 $D=0
M245 VSS 199 111 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=2945 $D=0
M246 111 199 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=3195 $D=0
M247 VSS 199 111 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=3445 $D=0
M248 112 200 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=3695 $D=0
M249 VSS 200 112 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=3945 $D=0
M250 112 200 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=4195 $D=0
M251 VSS 200 112 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=4445 $D=0
M252 113 201 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=4695 $D=0
M253 VSS 201 113 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=4945 $D=0
M254 113 201 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=5195 $D=0
M255 VSS 201 113 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=5445 $D=0
M256 114 202 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=5695 $D=0
M257 VSS 202 114 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=5945 $D=0
M258 114 202 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=6195 $D=0
M259 VSS 202 114 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=6445 $D=0
M260 115 203 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=6695 $D=0
M261 VSS 203 115 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=6945 $D=0
M262 115 203 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=7195 $D=0
M263 VSS 203 115 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=7445 $D=0
M264 116 204 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=7695 $D=0
M265 VSS 204 116 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=7945 $D=0
M266 116 204 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=8195 $D=0
M267 VSS 204 116 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=8445 $D=0
M268 125 205 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=8695 $D=0
M269 VSS 205 125 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=8945 $D=0
M270 125 205 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=9195 $D=0
M271 VSS 205 125 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=9445 $D=0
M272 126 206 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=9695 $D=0
M273 VSS 206 126 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=9945 $D=0
M274 126 206 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=10195 $D=0
M275 VSS 206 126 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=10445 $D=0
M276 127 207 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=10695 $D=0
M277 VSS 207 127 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=10945 $D=0
M278 127 207 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=11195 $D=0
M279 VSS 207 127 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=11445 $D=0
M280 128 208 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=11695 $D=0
M281 VSS 208 128 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=11945 $D=0
M282 128 208 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=12195 $D=0
M283 VSS 208 128 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=12445 $D=0
M284 129 209 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=12695 $D=0
M285 VSS 209 129 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=12945 $D=0
M286 129 209 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=13195 $D=0
M287 VSS 209 129 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=13445 $D=0
M288 130 210 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=13695 $D=0
M289 VSS 210 130 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=13945 $D=0
M290 130 210 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=14195 $D=0
M291 VSS 210 130 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=14445 $D=0
M292 131 211 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=14695 $D=0
M293 VSS 211 131 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=14945 $D=0
M294 131 211 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=15195 $D=0
M295 VSS 211 131 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=15445 $D=0
M296 132 212 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=15695 $D=0
M297 VSS 212 132 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=15945 $D=0
M298 132 212 VSS VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=16195 $D=0
M299 VSS 212 132 VSS n12ll L=6e-08 W=7.5e-07 $X=20700 $Y=16445 $D=0
M300 47 105 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=695 $D=0
M301 VSS 105 47 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=945 $D=0
M302 48 106 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=1195 $D=0
M303 VSS 106 48 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=1445 $D=0
M304 49 107 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=1695 $D=0
M305 VSS 107 49 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=1945 $D=0
M306 50 108 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=2195 $D=0
M307 VSS 108 50 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=2445 $D=0
M308 51 109 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=2695 $D=0
M309 VSS 109 51 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=2945 $D=0
M310 52 110 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=3195 $D=0
M311 VSS 110 52 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=3445 $D=0
M312 53 111 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=3695 $D=0
M313 VSS 111 53 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=3945 $D=0
M314 54 112 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=4195 $D=0
M315 VSS 112 54 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=4445 $D=0
M316 55 113 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=4695 $D=0
M317 VSS 113 55 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=4945 $D=0
M318 56 114 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=5195 $D=0
M319 VSS 114 56 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=5445 $D=0
M320 57 115 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=5695 $D=0
M321 VSS 115 57 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=5945 $D=0
M322 58 116 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=6195 $D=0
M323 VSS 116 58 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=6445 $D=0
M324 59 117 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=6695 $D=0
M325 VSS 117 59 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=6945 $D=0
M326 60 118 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=7195 $D=0
M327 VSS 118 60 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=7445 $D=0
M328 61 119 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=7695 $D=0
M329 VSS 119 61 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=7945 $D=0
M330 62 120 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=8195 $D=0
M331 VSS 120 62 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=8445 $D=0
M332 63 121 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=8695 $D=0
M333 VSS 121 63 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=8945 $D=0
M334 64 122 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=9195 $D=0
M335 VSS 122 64 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=9445 $D=0
M336 65 123 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=9695 $D=0
M337 VSS 123 65 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=9945 $D=0
M338 66 124 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=10195 $D=0
M339 VSS 124 66 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=10445 $D=0
M340 67 125 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=10695 $D=0
M341 VSS 125 67 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=10945 $D=0
M342 68 126 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=11195 $D=0
M343 VSS 126 68 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=11445 $D=0
M344 69 127 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=11695 $D=0
M345 VSS 127 69 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=11945 $D=0
M346 70 128 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=12195 $D=0
M347 VSS 128 70 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=12445 $D=0
M348 71 129 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=12695 $D=0
M349 VSS 129 71 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=12945 $D=0
M350 72 130 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=13195 $D=0
M351 VSS 130 72 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=13445 $D=0
M352 73 131 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=13695 $D=0
M353 VSS 131 73 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=13945 $D=0
M354 74 132 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=14195 $D=0
M355 VSS 132 74 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=14445 $D=0
M356 75 133 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=14695 $D=0
M357 VSS 133 75 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=14945 $D=0
M358 76 134 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=15195 $D=0
M359 VSS 134 76 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=15445 $D=0
M360 77 135 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=15695 $D=0
M361 VSS 135 77 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=15945 $D=0
M362 78 136 VSS VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=16195 $D=0
M363 VSS 136 78 VSS n12ll L=6e-08 W=1e-06 $X=22360 $Y=16445 $D=0
M364 2 105 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=695 $D=2
M365 VDD 105 2 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=945 $D=2
M366 3 106 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=1195 $D=2
M367 VDD 106 3 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=1445 $D=2
M368 4 107 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=1695 $D=2
M369 VDD 107 4 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=1945 $D=2
M370 5 108 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=2195 $D=2
M371 VDD 108 5 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=2445 $D=2
M372 6 109 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=2695 $D=2
M373 VDD 109 6 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=2945 $D=2
M374 7 110 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=3195 $D=2
M375 VDD 110 7 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=3445 $D=2
M376 8 111 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=3695 $D=2
M377 VDD 111 8 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=3945 $D=2
M378 9 112 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=4195 $D=2
M379 VDD 112 9 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=4445 $D=2
M380 10 113 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=4695 $D=2
M381 VDD 113 10 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=4945 $D=2
M382 11 114 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=5195 $D=2
M383 VDD 114 11 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=5445 $D=2
M384 12 115 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=5695 $D=2
M385 VDD 115 12 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=5945 $D=2
M386 13 116 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=6195 $D=2
M387 VDD 116 13 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=6445 $D=2
M388 14 117 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=6695 $D=2
M389 VDD 117 14 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=6945 $D=2
M390 15 118 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=7195 $D=2
M391 VDD 118 15 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=7445 $D=2
M392 16 119 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=7695 $D=2
M393 VDD 119 16 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=7945 $D=2
M394 17 120 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=8195 $D=2
M395 VDD 120 17 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=8445 $D=2
M396 18 121 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=8695 $D=2
M397 VDD 121 18 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=8945 $D=2
M398 19 122 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=9195 $D=2
M399 VDD 122 19 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=9445 $D=2
M400 20 123 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=9695 $D=2
M401 VDD 123 20 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=9945 $D=2
M402 21 124 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=10195 $D=2
M403 VDD 124 21 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=10445 $D=2
M404 22 125 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=10695 $D=2
M405 VDD 125 22 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=10945 $D=2
M406 23 126 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=11195 $D=2
M407 VDD 126 23 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=11445 $D=2
M408 24 127 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=11695 $D=2
M409 VDD 127 24 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=11945 $D=2
M410 25 128 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=12195 $D=2
M411 VDD 128 25 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=12445 $D=2
M412 26 129 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=12695 $D=2
M413 VDD 129 26 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=12945 $D=2
M414 27 130 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=13195 $D=2
M415 VDD 130 27 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=13445 $D=2
M416 28 131 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=13695 $D=2
M417 VDD 131 28 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=13945 $D=2
M418 29 132 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=14195 $D=2
M419 VDD 132 29 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=14445 $D=2
M420 30 133 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=14695 $D=2
M421 VDD 133 30 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=14945 $D=2
M422 31 134 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=15195 $D=2
M423 VDD 134 31 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=15445 $D=2
M424 32 135 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=15695 $D=2
M425 VDD 135 32 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=15945 $D=2
M426 33 136 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=16195 $D=2
M427 VDD 136 33 VDD p12ll L=6e-08 W=2.5e-06 $X=940 $Y=16445 $D=2
M428 105 137 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=695 $D=2
M429 VDD 137 105 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=945 $D=2
M430 105 137 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=1195 $D=2
M431 VDD 137 105 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=1445 $D=2
M432 106 138 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=1695 $D=2
M433 VDD 138 106 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=1945 $D=2
M434 106 138 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=2195 $D=2
M435 VDD 138 106 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=2445 $D=2
M436 107 139 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=2695 $D=2
M437 VDD 139 107 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=2945 $D=2
M438 107 139 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=3195 $D=2
M439 VDD 139 107 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=3445 $D=2
M440 108 140 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=3695 $D=2
M441 VDD 140 108 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=3945 $D=2
M442 108 140 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=4195 $D=2
M443 VDD 140 108 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=4445 $D=2
M444 117 141 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=4695 $D=2
M445 VDD 141 117 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=4945 $D=2
M446 117 141 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=5195 $D=2
M447 VDD 141 117 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=5445 $D=2
M448 118 142 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=5695 $D=2
M449 VDD 142 118 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=5945 $D=2
M450 118 142 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=6195 $D=2
M451 VDD 142 118 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=6445 $D=2
M452 119 143 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=6695 $D=2
M453 VDD 143 119 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=6945 $D=2
M454 119 143 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=7195 $D=2
M455 VDD 143 119 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=7445 $D=2
M456 120 144 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=7695 $D=2
M457 VDD 144 120 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=7945 $D=2
M458 120 144 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=8195 $D=2
M459 VDD 144 120 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=8445 $D=2
M460 121 145 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=8695 $D=2
M461 VDD 145 121 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=8945 $D=2
M462 121 145 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=9195 $D=2
M463 VDD 145 121 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=9445 $D=2
M464 122 146 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=9695 $D=2
M465 VDD 146 122 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=9945 $D=2
M466 122 146 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=10195 $D=2
M467 VDD 146 122 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=10445 $D=2
M468 123 147 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=10695 $D=2
M469 VDD 147 123 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=10945 $D=2
M470 123 147 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=11195 $D=2
M471 VDD 147 123 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=11445 $D=2
M472 124 148 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=11695 $D=2
M473 VDD 148 124 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=11945 $D=2
M474 124 148 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=12195 $D=2
M475 VDD 148 124 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=12445 $D=2
M476 133 149 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=12695 $D=2
M477 VDD 149 133 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=12945 $D=2
M478 133 149 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=13195 $D=2
M479 VDD 149 133 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=13445 $D=2
M480 134 150 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=13695 $D=2
M481 VDD 150 134 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=13945 $D=2
M482 134 150 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=14195 $D=2
M483 VDD 150 134 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=14445 $D=2
M484 135 151 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=14695 $D=2
M485 VDD 151 135 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=14945 $D=2
M486 135 151 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=15195 $D=2
M487 VDD 151 135 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=15445 $D=2
M488 136 152 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=15695 $D=2
M489 VDD 152 136 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=15945 $D=2
M490 136 152 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=16195 $D=2
M491 VDD 152 136 VDD p12ll L=6e-08 W=7.5e-07 $X=6950 $Y=16445 $D=2
M492 137 153 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=700 $D=2
M493 VDD 153 137 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=965 $D=2
M494 138 154 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=2175 $D=2
M495 VDD 154 138 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=2440 $D=2
M496 139 155 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=2700 $D=2
M497 VDD 155 139 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=2965 $D=2
M498 140 156 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=4175 $D=2
M499 VDD 156 140 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=4440 $D=2
M500 141 157 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=4700 $D=2
M501 VDD 157 141 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=4965 $D=2
M502 142 158 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=6175 $D=2
M503 VDD 158 142 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=6440 $D=2
M504 143 159 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=6700 $D=2
M505 VDD 159 143 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=6965 $D=2
M506 144 160 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=8175 $D=2
M507 VDD 160 144 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=8440 $D=2
M508 145 161 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=8700 $D=2
M509 VDD 161 145 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=8965 $D=2
M510 146 162 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=10175 $D=2
M511 VDD 162 146 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=10440 $D=2
M512 147 163 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=10700 $D=2
M513 VDD 163 147 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=10965 $D=2
M514 148 164 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=12175 $D=2
M515 VDD 164 148 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=12440 $D=2
M516 149 165 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=12700 $D=2
M517 VDD 165 149 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=12965 $D=2
M518 150 166 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=14175 $D=2
M519 VDD 166 150 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=14440 $D=2
M520 151 167 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=14700 $D=2
M521 VDD 167 151 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=14965 $D=2
M522 152 168 VDD VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=16175 $D=2
M523 VDD 168 152 VDD p12ll L=6e-08 W=4e-07 $X=8220 $Y=16440 $D=2
M524 153 177 35 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=1180 $D=2
M525 VDD 173 153 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=1440 $D=2
M526 154 173 VDD VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=1700 $D=2
M527 36 177 154 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=1960 $D=2
M528 155 177 37 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=3180 $D=2
M529 VDD 173 155 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=3440 $D=2
M530 156 173 VDD VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=3700 $D=2
M531 38 177 156 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=3960 $D=2
M532 157 178 38 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=5180 $D=2
M533 VDD 174 157 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=5440 $D=2
M534 158 174 VDD VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=5700 $D=2
M535 37 178 158 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=5960 $D=2
M536 159 178 36 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=7180 $D=2
M537 VDD 174 159 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=7440 $D=2
M538 160 174 VDD VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=7700 $D=2
M539 35 178 160 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=7960 $D=2
M540 161 179 35 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=9180 $D=2
M541 VDD 175 161 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=9440 $D=2
M542 162 175 VDD VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=9700 $D=2
M543 36 179 162 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=9960 $D=2
M544 163 179 37 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=11180 $D=2
M545 VDD 175 163 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=11440 $D=2
M546 164 175 VDD VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=11700 $D=2
M547 38 179 164 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=11960 $D=2
M548 165 180 38 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=13180 $D=2
M549 VDD 176 165 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=13440 $D=2
M550 166 176 VDD VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=13700 $D=2
M551 37 180 166 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=13960 $D=2
M552 167 180 36 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=15180 $D=2
M553 VDD 176 167 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=15440 $D=2
M554 168 176 VDD VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=15700 $D=2
M555 35 180 168 VDD p12ll L=6e-08 W=4e-07 $X=8960 $Y=15960 $D=2
M556 177 173 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=1120 $D=2
M557 VDD 173 177 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=1405 $D=2
M558 177 173 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=1695 $D=2
M559 VDD 173 177 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=1985 $D=2
M560 173 169 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=2275 $D=2
M561 VDD 169 173 VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=2560 $D=2
M562 173 169 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=2850 $D=2
M563 VDD 169 173 VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=3140 $D=2
M564 169 39 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=3430 $D=2
M565 VDD 40 169 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=3720 $D=2
M566 169 VDD VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=4010 $D=2
M567 VDD VDD 170 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=5130 $D=2
M568 170 40 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=5420 $D=2
M569 VDD 41 170 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=5710 $D=2
M570 174 170 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=6000 $D=2
M571 VDD 170 174 VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=6290 $D=2
M572 174 170 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=6580 $D=2
M573 VDD 170 174 VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=6865 $D=2
M574 178 174 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=7155 $D=2
M575 VDD 174 178 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=7445 $D=2
M576 178 174 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=7735 $D=2
M577 VDD 174 178 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=8020 $D=2
M578 179 175 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=9120 $D=2
M579 VDD 175 179 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=9405 $D=2
M580 179 175 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=9695 $D=2
M581 VDD 175 179 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=9985 $D=2
M582 175 171 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=10275 $D=2
M583 VDD 171 175 VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=10560 $D=2
M584 175 171 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=10850 $D=2
M585 VDD 171 175 VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=11140 $D=2
M586 171 39 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=11430 $D=2
M587 VDD 42 171 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=11720 $D=2
M588 171 VDD VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=12010 $D=2
M589 VDD VDD 172 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=13130 $D=2
M590 172 42 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=13420 $D=2
M591 VDD 41 172 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=13710 $D=2
M592 176 172 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=14000 $D=2
M593 VDD 172 176 VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=14290 $D=2
M594 176 172 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=14580 $D=2
M595 VDD 172 176 VDD p12ll L=6e-08 W=7.5e-07 $X=14015 $Y=14865 $D=2
M596 180 176 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=15155 $D=2
M597 VDD 176 180 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=15445 $D=2
M598 180 176 VDD VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=15735 $D=2
M599 VDD 176 180 VDD p12ll L=6e-08 W=5e-07 $X=14015 $Y=16020 $D=2
M600 181 177 43 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=1180 $D=2
M601 VDD 173 181 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=1440 $D=2
M602 182 173 VDD VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=1700 $D=2
M603 44 177 182 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=1960 $D=2
M604 183 177 45 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=3180 $D=2
M605 VDD 173 183 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=3440 $D=2
M606 184 173 VDD VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=3700 $D=2
M607 46 177 184 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=3960 $D=2
M608 185 178 46 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=5180 $D=2
M609 VDD 174 185 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=5440 $D=2
M610 186 174 VDD VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=5700 $D=2
M611 45 178 186 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=5960 $D=2
M612 187 178 44 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=7180 $D=2
M613 VDD 174 187 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=7440 $D=2
M614 188 174 VDD VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=7700 $D=2
M615 43 178 188 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=7960 $D=2
M616 189 179 43 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=9180 $D=2
M617 VDD 175 189 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=9440 $D=2
M618 190 175 VDD VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=9700 $D=2
M619 44 179 190 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=9960 $D=2
M620 191 179 45 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=11180 $D=2
M621 VDD 175 191 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=11440 $D=2
M622 192 175 VDD VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=11700 $D=2
M623 46 179 192 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=11960 $D=2
M624 193 180 46 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=13180 $D=2
M625 VDD 176 193 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=13440 $D=2
M626 194 176 VDD VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=13700 $D=2
M627 45 180 194 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=13960 $D=2
M628 195 180 44 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=15180 $D=2
M629 VDD 176 195 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=15440 $D=2
M630 196 176 VDD VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=15700 $D=2
M631 43 180 196 VDD p12ll L=6e-08 W=4e-07 $X=17890 $Y=15960 $D=2
M632 197 181 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=700 $D=2
M633 VDD 181 197 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=965 $D=2
M634 198 182 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=2175 $D=2
M635 VDD 182 198 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=2440 $D=2
M636 199 183 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=2700 $D=2
M637 VDD 183 199 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=2965 $D=2
M638 200 184 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=4175 $D=2
M639 VDD 184 200 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=4440 $D=2
M640 201 185 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=4700 $D=2
M641 VDD 185 201 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=4965 $D=2
M642 202 186 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=6175 $D=2
M643 VDD 186 202 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=6440 $D=2
M644 203 187 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=6700 $D=2
M645 VDD 187 203 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=6965 $D=2
M646 204 188 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=8175 $D=2
M647 VDD 188 204 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=8440 $D=2
M648 205 189 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=8700 $D=2
M649 VDD 189 205 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=8965 $D=2
M650 206 190 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=10175 $D=2
M651 VDD 190 206 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=10440 $D=2
M652 207 191 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=10700 $D=2
M653 VDD 191 207 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=10965 $D=2
M654 208 192 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=12175 $D=2
M655 VDD 192 208 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=12440 $D=2
M656 209 193 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=12700 $D=2
M657 VDD 193 209 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=12965 $D=2
M658 210 194 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=14175 $D=2
M659 VDD 194 210 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=14440 $D=2
M660 211 195 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=14700 $D=2
M661 VDD 195 211 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=14965 $D=2
M662 212 196 VDD VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=16175 $D=2
M663 VDD 196 212 VDD p12ll L=6e-08 W=4e-07 $X=18630 $Y=16440 $D=2
M664 109 197 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=695 $D=2
M665 VDD 197 109 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=945 $D=2
M666 109 197 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=1195 $D=2
M667 VDD 197 109 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=1445 $D=2
M668 110 198 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=1695 $D=2
M669 VDD 198 110 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=1945 $D=2
M670 110 198 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=2195 $D=2
M671 VDD 198 110 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=2445 $D=2
M672 111 199 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=2695 $D=2
M673 VDD 199 111 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=2945 $D=2
M674 111 199 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=3195 $D=2
M675 VDD 199 111 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=3445 $D=2
M676 112 200 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=3695 $D=2
M677 VDD 200 112 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=3945 $D=2
M678 112 200 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=4195 $D=2
M679 VDD 200 112 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=4445 $D=2
M680 113 201 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=4695 $D=2
M681 VDD 201 113 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=4945 $D=2
M682 113 201 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=5195 $D=2
M683 VDD 201 113 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=5445 $D=2
M684 114 202 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=5695 $D=2
M685 VDD 202 114 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=5945 $D=2
M686 114 202 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=6195 $D=2
M687 VDD 202 114 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=6445 $D=2
M688 115 203 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=6695 $D=2
M689 VDD 203 115 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=6945 $D=2
M690 115 203 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=7195 $D=2
M691 VDD 203 115 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=7445 $D=2
M692 116 204 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=7695 $D=2
M693 VDD 204 116 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=7945 $D=2
M694 116 204 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=8195 $D=2
M695 VDD 204 116 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=8445 $D=2
M696 125 205 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=8695 $D=2
M697 VDD 205 125 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=8945 $D=2
M698 125 205 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=9195 $D=2
M699 VDD 205 125 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=9445 $D=2
M700 126 206 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=9695 $D=2
M701 VDD 206 126 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=9945 $D=2
M702 126 206 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=10195 $D=2
M703 VDD 206 126 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=10445 $D=2
M704 127 207 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=10695 $D=2
M705 VDD 207 127 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=10945 $D=2
M706 127 207 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=11195 $D=2
M707 VDD 207 127 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=11445 $D=2
M708 128 208 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=11695 $D=2
M709 VDD 208 128 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=11945 $D=2
M710 128 208 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=12195 $D=2
M711 VDD 208 128 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=12445 $D=2
M712 129 209 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=12695 $D=2
M713 VDD 209 129 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=12945 $D=2
M714 129 209 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=13195 $D=2
M715 VDD 209 129 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=13445 $D=2
M716 130 210 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=13695 $D=2
M717 VDD 210 130 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=13945 $D=2
M718 130 210 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=14195 $D=2
M719 VDD 210 130 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=14445 $D=2
M720 131 211 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=14695 $D=2
M721 VDD 211 131 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=14945 $D=2
M722 131 211 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=15195 $D=2
M723 VDD 211 131 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=15445 $D=2
M724 132 212 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=15695 $D=2
M725 VDD 212 132 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=15945 $D=2
M726 132 212 VDD VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=16195 $D=2
M727 VDD 212 132 VDD p12ll L=6e-08 W=7.5e-07 $X=19550 $Y=16445 $D=2
M728 47 105 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=695 $D=2
M729 VDD 105 47 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=945 $D=2
M730 48 106 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=1195 $D=2
M731 VDD 106 48 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=1445 $D=2
M732 49 107 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=1695 $D=2
M733 VDD 107 49 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=1945 $D=2
M734 50 108 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=2195 $D=2
M735 VDD 108 50 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=2445 $D=2
M736 51 109 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=2695 $D=2
M737 VDD 109 51 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=2945 $D=2
M738 52 110 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=3195 $D=2
M739 VDD 110 52 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=3445 $D=2
M740 53 111 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=3695 $D=2
M741 VDD 111 53 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=3945 $D=2
M742 54 112 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=4195 $D=2
M743 VDD 112 54 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=4445 $D=2
M744 55 113 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=4695 $D=2
M745 VDD 113 55 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=4945 $D=2
M746 56 114 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=5195 $D=2
M747 VDD 114 56 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=5445 $D=2
M748 57 115 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=5695 $D=2
M749 VDD 115 57 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=5945 $D=2
M750 58 116 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=6195 $D=2
M751 VDD 116 58 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=6445 $D=2
M752 59 117 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=6695 $D=2
M753 VDD 117 59 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=6945 $D=2
M754 60 118 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=7195 $D=2
M755 VDD 118 60 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=7445 $D=2
M756 61 119 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=7695 $D=2
M757 VDD 119 61 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=7945 $D=2
M758 62 120 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=8195 $D=2
M759 VDD 120 62 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=8445 $D=2
M760 63 121 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=8695 $D=2
M761 VDD 121 63 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=8945 $D=2
M762 64 122 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=9195 $D=2
M763 VDD 122 64 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=9445 $D=2
M764 65 123 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=9695 $D=2
M765 VDD 123 65 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=9945 $D=2
M766 66 124 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=10195 $D=2
M767 VDD 124 66 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=10445 $D=2
M768 67 125 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=10695 $D=2
M769 VDD 125 67 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=10945 $D=2
M770 68 126 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=11195 $D=2
M771 VDD 126 68 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=11445 $D=2
M772 69 127 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=11695 $D=2
M773 VDD 127 69 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=11945 $D=2
M774 70 128 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=12195 $D=2
M775 VDD 128 70 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=12445 $D=2
M776 71 129 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=12695 $D=2
M777 VDD 129 71 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=12945 $D=2
M778 72 130 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=13195 $D=2
M779 VDD 130 72 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=13445 $D=2
M780 73 131 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=13695 $D=2
M781 VDD 131 73 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=13945 $D=2
M782 74 132 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=14195 $D=2
M783 VDD 132 74 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=14445 $D=2
M784 75 133 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=14695 $D=2
M785 VDD 133 75 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=14945 $D=2
M786 76 134 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=15195 $D=2
M787 VDD 134 76 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=15445 $D=2
M788 77 135 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=15695 $D=2
M789 VDD 135 77 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=15945 $D=2
M790 78 136 VDD VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=16195 $D=2
M791 VDD 136 78 VDD p12ll L=6e-08 W=2.5e-06 $X=23810 $Y=16445 $D=2
.ENDS
***************************************
.SUBCKT XDEC64_VHSSP 1 2 3 4 5 6 7 8 9 10 11 12 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43
+ 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147
** N=166 EP=144 IP=208 FDC=1584
X0 7 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38
+ 39 40 41 42 43 44 45 46 47 48 49 50 51 8 11 12 10 9 1 5
+ 2 6 17 18 16 19 52 53 54 55 56 57 58 59 60 61 62 63 64 65
+ 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ LEAF_XDEC4_VHSSRAM $T=0 0 0 0 $X=-1400 $Y=-350
X1 7 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 8 11 12 10 9 1 4
+ 2 3 17 18 16 19 116 117 118 119 120 121 122 123 124 125 126 127 128 129
+ 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147
+ LEAF_XDEC4_VHSSRAM $T=0 17200 0 0 $X=-1400 $Y=16850
.ENDS
***************************************
.SUBCKT SOP_DC_X128Y8_620 VSS VDD 5 13 EMCLK
** N=100 EP=5 IP=0 FDC=140
*.CALIBRE ISOLATED NETS: A[8] A[9] A[6] A[7] A[3] A[4] A[5] CEN CLK A[2] A[0] A[1] WEN
M0 5 21 VSS VSS n12ll L=6e-08 W=1e-06 $X=3730 $Y=1665 $D=0
M1 VSS 30 28 VSS n12ll L=6e-08 W=5e-07 $X=6195 $Y=2390 $D=0
M2 28 30 VSS VSS n12ll L=6e-08 W=5e-07 $X=6195 $Y=2680 $D=0
M3 VSS 30 28 VSS n12ll L=6e-08 W=5e-07 $X=6195 $Y=2980 $D=0
M4 29 29 VSS VSS n12ll L=6e-08 W=5e-07 $X=6195 $Y=3270 $D=0
M5 VSS 29 29 VSS n12ll L=6e-08 W=5e-07 $X=6195 $Y=3570 $D=0
M6 VSS 28 32 VSS n12ll L=6e-08 W=4e-07 $X=10080 $Y=2135 $D=0
M7 33 32 VSS VSS n12ll L=6e-08 W=4e-07 $X=10370 $Y=2135 $D=0
M8 VSS 28 35 VSS n12ll L=6e-08 W=4e-07 $X=12560 $Y=2165 $D=0
M9 37 35 VSS VSS n12ll L=6e-08 W=4e-07 $X=12850 $Y=2165 $D=0
M10 85 32 39 VSS n12ll L=6e-08 W=4e-07 $X=13445 $Y=2150 $D=0
M11 86 50 85 VSS n12ll L=6e-08 W=4e-07 $X=13735 $Y=2150 $D=0
M12 VSS 35 86 VSS n12ll L=6e-08 W=4e-07 $X=14025 $Y=2150 $D=0
M13 87 35 VSS VSS n12ll L=6e-08 W=4e-07 $X=14320 $Y=2150 $D=0
M14 40 50 87 VSS n12ll L=6e-08 W=4e-07 $X=14610 $Y=2150 $D=0
M15 88 50 42 VSS n12ll L=6e-08 W=4e-07 $X=15240 $Y=2090 $D=0
M16 VSS 43 88 VSS n12ll L=6e-08 W=4e-07 $X=15530 $Y=2090 $D=0
M17 89 33 VSS VSS n12ll L=6e-08 W=4e-07 $X=15830 $Y=2090 $D=0
M18 43 37 89 VSS n12ll L=6e-08 W=4e-07 $X=16120 $Y=2090 $D=0
M19 45 37 VSS VSS n12ll L=6e-08 W=4e-07 $X=16750 $Y=2090 $D=0
M20 VSS 33 45 VSS n12ll L=6e-08 W=4e-07 $X=17040 $Y=2090 $D=0
M21 46 45 VSS VSS n12ll L=6e-08 W=4e-07 $X=17340 $Y=2090 $D=0
M22 VSS 50 46 VSS n12ll L=6e-08 W=4e-07 $X=17630 $Y=2090 $D=0
M23 48 35 VSS VSS n12ll L=6e-08 W=4e-07 $X=18260 $Y=2150 $D=0
M24 VSS 50 48 VSS n12ll L=6e-08 W=4e-07 $X=18550 $Y=2150 $D=0
M25 VSS 50 49 VSS n12ll L=6e-08 W=4e-07 $X=19235 $Y=2115 $D=0
M26 50 28 VSS VSS n12ll L=6e-08 W=4e-07 $X=19525 $Y=2115 $D=0
M27 34 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=12055 $Y=3515 $D=96
M28 34 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=12055 $Y=3840 $D=96
M29 34 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=12055 $Y=4305 $D=96
M30 34 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=12055 $Y=4630 $D=96
M31 13 EMCLK 36 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=13160 $Y=3515 $D=96
M32 13 EMCLK 36 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=13160 $Y=3840 $D=96
M33 13 EMCLK 36 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=13160 $Y=4305 $D=96
M34 13 EMCLK 36 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=13160 $Y=4630 $D=96
M35 38 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=13535 $Y=3515 $D=96
M36 38 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=13535 $Y=3840 $D=96
M37 38 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=13535 $Y=4305 $D=96
M38 38 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=13535 $Y=4630 $D=96
M39 13 EMCLK 41 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=14640 $Y=3515 $D=96
M40 13 EMCLK 41 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=14640 $Y=3840 $D=96
M41 13 EMCLK 41 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=14640 $Y=4305 $D=96
M42 13 EMCLK 41 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=14640 $Y=4630 $D=96
M43 41 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=15015 $Y=3515 $D=96
M44 41 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=15015 $Y=3840 $D=96
M45 41 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=15015 $Y=4305 $D=96
M46 41 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=15015 $Y=4630 $D=96
M47 13 EMCLK 44 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=16120 $Y=3515 $D=96
M48 13 EMCLK 44 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=16120 $Y=3840 $D=96
M49 13 EMCLK 44 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=16120 $Y=4305 $D=96
M50 13 EMCLK 44 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=16120 $Y=4630 $D=96
M51 44 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=16495 $Y=3515 $D=96
M52 44 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=16495 $Y=3840 $D=96
M53 44 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=16495 $Y=4305 $D=96
M54 44 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=16495 $Y=4630 $D=96
M55 13 EMCLK 47 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=17600 $Y=3515 $D=96
M56 13 EMCLK 47 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=17600 $Y=3840 $D=96
M57 13 EMCLK 47 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=17600 $Y=4305 $D=96
M58 13 EMCLK 47 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=17600 $Y=4630 $D=96
M59 47 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=17975 $Y=3515 $D=96
M60 47 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=17975 $Y=3840 $D=96
M61 47 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=17975 $Y=4305 $D=96
M62 47 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=17975 $Y=4630 $D=96
M63 13 EMCLK 51 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=19080 $Y=3515 $D=96
M64 13 EMCLK 51 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=19080 $Y=3840 $D=96
M65 13 EMCLK 51 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=19080 $Y=4305 $D=96
M66 13 EMCLK 51 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=19080 $Y=4630 $D=96
M67 51 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=19455 $Y=3515 $D=96
M68 51 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=19455 $Y=3840 $D=96
M69 51 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=19455 $Y=4305 $D=96
M70 51 EMCLK 13 VSS DNNPGSVT L=7.5e-08 W=1.25e-07 $X=19455 $Y=4630 $D=96
M71 VSS VDD 34 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=12420 $Y=3430 $D=95
M72 VSS VDD 34 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=12420 $Y=3840 $D=95
M73 VSS VDD 34 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=12420 $Y=4220 $D=95
M74 VSS VDD 34 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=12420 $Y=4630 $D=95
M75 36 39 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=12805 $Y=3430 $D=95
M76 36 39 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=12805 $Y=3840 $D=95
M77 36 39 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=12805 $Y=4220 $D=95
M78 36 39 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=12805 $Y=4630 $D=95
M79 VSS 40 38 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=13900 $Y=3430 $D=95
M80 VSS 40 38 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=13900 $Y=3840 $D=95
M81 VSS 40 38 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=13900 $Y=4220 $D=95
M82 VSS 40 38 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=13900 $Y=4630 $D=95
M83 41 42 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=14285 $Y=3430 $D=95
M84 41 42 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=14285 $Y=3840 $D=95
M85 41 42 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=14285 $Y=4220 $D=95
M86 41 42 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=14285 $Y=4630 $D=95
M87 VSS 42 41 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=15380 $Y=3430 $D=95
M88 VSS 42 41 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=15380 $Y=3840 $D=95
M89 VSS 42 41 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=15380 $Y=4220 $D=95
M90 VSS 42 41 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=15380 $Y=4630 $D=95
M91 44 46 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=15765 $Y=3430 $D=95
M92 44 46 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=15765 $Y=3840 $D=95
M93 44 46 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=15765 $Y=4220 $D=95
M94 44 46 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=15765 $Y=4630 $D=95
M95 VSS 46 44 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=16860 $Y=3430 $D=95
M96 VSS 46 44 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=16860 $Y=3840 $D=95
M97 VSS 46 44 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=16860 $Y=4220 $D=95
M98 VSS 46 44 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=16860 $Y=4630 $D=95
M99 47 48 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=17245 $Y=3430 $D=95
M100 47 48 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=17245 $Y=3840 $D=95
M101 47 48 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=17245 $Y=4220 $D=95
M102 47 48 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=17245 $Y=4630 $D=95
M103 VSS 48 47 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=18340 $Y=3430 $D=95
M104 VSS 48 47 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=18340 $Y=3840 $D=95
M105 VSS 48 47 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=18340 $Y=4220 $D=95
M106 VSS 48 47 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=18340 $Y=4630 $D=95
M107 51 49 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=18725 $Y=3430 $D=95
M108 51 49 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=18725 $Y=3840 $D=95
M109 51 49 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=18725 $Y=4220 $D=95
M110 51 49 VSS VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=18725 $Y=4630 $D=95
M111 VSS 49 51 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=19820 $Y=3430 $D=95
M112 VSS 49 51 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=19820 $Y=3840 $D=95
M113 VSS 49 51 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=19820 $Y=4220 $D=95
M114 VSS 49 51 VSS DNNPDSVT L=6.5e-08 W=2.1e-07 $X=19820 $Y=4630 $D=95
M115 21 21 VDD VDD p12ll L=6e-08 W=4e-07 $X=2560 $Y=1665 $D=2
M116 VDD 30 30 VDD p12ll L=6e-08 W=1e-06 $X=7495 $Y=2980 $D=2
M117 31 29 VDD VDD p12ll L=6e-08 W=1e-06 $X=7495 $Y=3270 $D=2
M118 VDD 29 31 VDD p12ll L=6e-08 W=1e-06 $X=7495 $Y=3570 $D=2
M119 VDD 28 32 VDD p12ll L=6e-08 W=4e-07 $X=10080 $Y=1240 $D=2
M120 33 32 VDD VDD p12ll L=6e-08 W=4e-07 $X=10370 $Y=1240 $D=2
M121 VDD 28 35 VDD p12ll L=6e-08 W=4e-07 $X=12560 $Y=1055 $D=2
M122 37 35 VDD VDD p12ll L=6e-08 W=4e-07 $X=12850 $Y=1055 $D=2
M123 VDD 32 39 VDD p12ll L=6e-08 W=4e-07 $X=13445 $Y=1070 $D=2
M124 39 50 VDD VDD p12ll L=6e-08 W=4e-07 $X=13735 $Y=1070 $D=2
M125 VDD 35 39 VDD p12ll L=6e-08 W=4e-07 $X=14025 $Y=1070 $D=2
M126 40 35 VDD VDD p12ll L=6e-08 W=4e-07 $X=14320 $Y=1070 $D=2
M127 VDD 50 40 VDD p12ll L=6e-08 W=4e-07 $X=14610 $Y=1070 $D=2
M128 42 50 VDD VDD p12ll L=6e-08 W=4e-07 $X=15240 $Y=1040 $D=2
M129 VDD 43 42 VDD p12ll L=6e-08 W=4e-07 $X=15530 $Y=1040 $D=2
M130 43 33 VDD VDD p12ll L=6e-08 W=4e-07 $X=15830 $Y=1040 $D=2
M131 VDD 37 43 VDD p12ll L=6e-08 W=4e-07 $X=16120 $Y=1040 $D=2
M132 98 37 45 VDD p12ll L=6e-08 W=4e-07 $X=16750 $Y=1040 $D=2
M133 VDD 33 98 VDD p12ll L=6e-08 W=4e-07 $X=17040 $Y=1040 $D=2
M134 99 45 VDD VDD p12ll L=6e-08 W=4e-07 $X=17340 $Y=1040 $D=2
M135 46 50 99 VDD p12ll L=6e-08 W=4e-07 $X=17630 $Y=1040 $D=2
M136 100 35 48 VDD p12ll L=6e-08 W=4e-07 $X=18260 $Y=1040 $D=2
M137 VDD 50 100 VDD p12ll L=6e-08 W=4e-07 $X=18550 $Y=1040 $D=2
M138 VDD 50 49 VDD p12ll L=6e-08 W=4e-07 $X=19235 $Y=1035 $D=2
M139 50 28 VDD VDD p12ll L=6e-08 W=4e-07 $X=19525 $Y=1035 $D=2
.ENDS
***************************************
.SUBCKT Logic_leafcell_X128Y8_VHS vdd vss RDE PXB[3] A[8] PXB[2] PXB[1] PXB[0] A[9] A[6] PXA[3] PXA[2] PXA[1] PXA[0] A[7] FCKX[3] ZASX ZAS FCKX[2] A[5]
+ A[3] CEN FCKX[0] CLK FCKX[1] EMCLK DBL FCKX[7] FCKX[6] FCKX[4] FCKX[5] A[4] YX[3] DCTRCLK RWLL YX[2] WEN DCTRCLKX SACK4 YX[0]
+ YX[1] A[2] SACK1 YX[7] A[0] YX[6] WE A[1] YX[4] RWLR YX[5]
** N=436 EP=51 IP=0 FDC=985
M0 343 vdd vss vss n12ll L=3e-07 W=4e-07 $X=610 $Y=2925 $D=0
M1 124 126 vss vss n12ll L=6e-07 W=1.2e-07 $X=1100 $Y=3835 $D=0
M2 99 RDE 343 vss n12ll L=6e-08 W=4e-07 $X=1110 $Y=2925 $D=0
M3 114 99 vss vss n12ll L=6e-08 W=4e-07 $X=1700 $Y=2940 $D=0
M4 vss 114 115 vss n12ll L=6e-08 W=4e-07 $X=2320 $Y=2940 $D=0
M5 PXB[3] 118 vss vss n12ll L=6e-08 W=1.5e-06 $X=2590 $Y=24740 $D=0
M6 119 115 vss vss n12ll L=6e-08 W=4e-07 $X=2600 $Y=2940 $D=0
M7 123 PXB[2] vss vss n12ll L=6e-07 W=1.2e-07 $X=2670 $Y=23955 $D=0
M8 353 135 116 vss n12ll L=6e-08 W=1.495e-06 $X=2710 $Y=12950 $D=0
M9 354 A[8] 117 vss n12ll L=6e-08 W=4e-07 $X=2730 $Y=7240 $D=0
M10 118 121 116 vss n12ll L=6e-08 W=2.5e-06 $X=2735 $Y=17190 $D=0
M11 vss PXB[3] 118 vss n12ll L=6e-07 W=1.2e-07 $X=2840 $Y=23305 $D=0
M12 vss 118 PXB[3] vss n12ll L=6e-08 W=1.5e-06 $X=2880 $Y=24740 $D=0
M13 vss 130 353 vss n12ll L=6e-08 W=1.495e-06 $X=2890 $Y=12950 $D=0
M14 vss 117 135 vss n12ll L=6e-08 W=7e-07 $X=2925 $Y=11400 $D=0
M15 vss vss A[8] vss n12ll L=6e-08 W=2e-07 $X=2935 $Y=5860 $D=0
M16 vss vdd 354 vss n12ll L=3e-07 W=4e-07 $X=3045 $Y=7240 $D=0
M17 124 121 119 vss n12ll L=6e-08 W=1e-06 $X=3060 $Y=2690 $D=0
M18 355 130 vss vss n12ll L=6e-08 W=1.495e-06 $X=3160 $Y=12950 $D=0
M19 PXB[2] 123 vss vss n12ll L=6e-08 W=1.5e-06 $X=3170 $Y=24740 $D=0
M20 125 135 vss vss n12ll L=6e-08 W=7e-07 $X=3215 $Y=11400 $D=0
M21 122 121 123 vss n12ll L=6e-08 W=2.5e-06 $X=3315 $Y=17190 $D=0
M22 122 125 355 vss n12ll L=6e-08 W=1.495e-06 $X=3340 $Y=12950 $D=0
M23 vss 123 PXB[2] vss n12ll L=6e-08 W=1.5e-06 $X=3460 $Y=24740 $D=0
M24 vss 124 126 vss n12ll L=6e-08 W=4e-07 $X=3670 $Y=3120 $D=0
M25 PXB[0] 127 vss vss n12ll L=6e-08 W=1.5e-06 $X=3800 $Y=24740 $D=0
M26 132 PXB[1] vss vss n12ll L=6e-07 W=1.2e-07 $X=3880 $Y=23305 $D=0
M27 356 125 128 vss n12ll L=6e-08 W=1.495e-06 $X=3920 $Y=12950 $D=0
M28 127 121 128 vss n12ll L=6e-08 W=2.5e-06 $X=3945 $Y=17190 $D=0
M29 129 126 vss vss n12ll L=6e-08 W=4e-07 $X=3950 $Y=3120 $D=0
M30 357 vdd vss vss n12ll L=3e-07 W=4e-07 $X=3995 $Y=7240 $D=0
M31 vss 133 130 vss n12ll L=6e-08 W=7e-07 $X=4045 $Y=11400 $D=0
M32 vss PXB[0] 127 vss n12ll L=6e-07 W=1.2e-07 $X=4050 $Y=23955 $D=0
M33 vss 127 PXB[0] vss n12ll L=6e-08 W=1.5e-06 $X=4090 $Y=24740 $D=0
M34 vss 131 356 vss n12ll L=6e-08 W=1.495e-06 $X=4100 $Y=12950 $D=0
M35 131 130 vss vss n12ll L=6e-08 W=7e-07 $X=4335 $Y=11400 $D=0
M36 358 131 vss vss n12ll L=6e-08 W=1.495e-06 $X=4370 $Y=12950 $D=0
M37 PXB[1] 132 vss vss n12ll L=6e-08 W=1.5e-06 $X=4380 $Y=24740 $D=0
M38 134 121 132 vss n12ll L=6e-08 W=2.5e-06 $X=4525 $Y=17190 $D=0
M39 133 A[9] 357 vss n12ll L=6e-08 W=4e-07 $X=4550 $Y=7240 $D=0
M40 134 135 358 vss n12ll L=6e-08 W=1.495e-06 $X=4550 $Y=12950 $D=0
M41 vss 132 PXB[1] vss n12ll L=6e-08 W=1.5e-06 $X=4670 $Y=24740 $D=0
M42 vss vss A[9] vss n12ll L=6e-08 W=2e-07 $X=4870 $Y=5860 $D=0
M43 vss A[6] 137 vss n12ll L=6e-08 W=4e-07 $X=4975 $Y=2655 $D=0
M44 PXA[3] 139 vss vss n12ll L=6e-08 W=1.5e-06 $X=5010 $Y=24740 $D=0
M45 142 PXA[2] vss vss n12ll L=6e-07 W=1.2e-07 $X=5090 $Y=23955 $D=0
M46 359 152 138 vss n12ll L=6e-08 W=1.495e-06 $X=5130 $Y=12950 $D=0
M47 139 121 138 vss n12ll L=6e-08 W=2.5e-06 $X=5155 $Y=17190 $D=0
M48 152 140 vss vss n12ll L=6e-08 W=5e-07 $X=5165 $Y=11400 $D=0
M49 vss PXA[3] 139 vss n12ll L=6e-07 W=1.2e-07 $X=5260 $Y=23300 $D=0
M50 vss 139 PXA[3] vss n12ll L=6e-08 W=1.5e-06 $X=5300 $Y=24740 $D=0
M51 vss 150 359 vss n12ll L=6e-08 W=1.495e-06 $X=5310 $Y=12950 $D=0
M52 145 137 vss vss n12ll L=3e-07 W=4e-07 $X=5335 $Y=2655 $D=0
M53 vss A[6] 140 vss n12ll L=6e-08 W=4e-07 $X=5375 $Y=7215 $D=0
M54 vss RDE 152 vss n12ll L=6e-08 W=5e-07 $X=5455 $Y=11400 $D=0
M55 360 150 vss vss n12ll L=6e-08 W=1.495e-06 $X=5580 $Y=12950 $D=0
M56 PXA[2] 142 vss vss n12ll L=6e-08 W=1.5e-06 $X=5590 $Y=24740 $D=0
M57 143 140 vss vss n12ll L=6e-08 W=4e-07 $X=5655 $Y=7215 $D=0
M58 141 121 142 vss n12ll L=6e-08 W=2.5e-06 $X=5735 $Y=17190 $D=0
M59 144 RDE vss vss n12ll L=6e-08 W=7e-07 $X=5745 $Y=11400 $D=0
M60 141 144 360 vss n12ll L=6e-08 W=1.495e-06 $X=5760 $Y=12950 $D=0
M61 vss vss A[6] vss n12ll L=6e-08 W=2e-07 $X=5810 $Y=5860 $D=0
M62 vss 142 PXA[2] vss n12ll L=6e-08 W=1.5e-06 $X=5880 $Y=24740 $D=0
M63 vss 143 144 vss n12ll L=6e-08 W=7e-07 $X=6035 $Y=11400 $D=0
M64 A[7] vss vss vss n12ll L=6e-08 W=2e-07 $X=6090 $Y=5860 $D=0
M65 PXA[0] 146 vss vss n12ll L=6e-08 W=1.5e-06 $X=6220 $Y=24740 $D=0
M66 148 145 vss vss n12ll L=6e-08 W=4e-07 $X=6285 $Y=2650 $D=0
M67 149 PXA[1] vss vss n12ll L=6e-07 W=1.2e-07 $X=6300 $Y=23300 $D=0
M68 361 144 147 vss n12ll L=6e-08 W=1.495e-06 $X=6340 $Y=12950 $D=0
M69 146 121 147 vss n12ll L=6e-08 W=2.5e-06 $X=6365 $Y=17190 $D=0
M70 362 vdd vss vss n12ll L=3e-07 W=4e-07 $X=6425 $Y=7215 $D=0
M71 vss PXA[0] 146 vss n12ll L=6e-07 W=1.2e-07 $X=6470 $Y=23955 $D=0
M72 vss 146 PXA[0] vss n12ll L=6e-08 W=1.5e-06 $X=6510 $Y=24740 $D=0
M73 vss 154 361 vss n12ll L=6e-08 W=1.495e-06 $X=6520 $Y=12950 $D=0
M74 363 154 vss vss n12ll L=6e-08 W=1.495e-06 $X=6790 $Y=12950 $D=0
M75 PXA[1] 149 vss vss n12ll L=6e-08 W=1.5e-06 $X=6800 $Y=24740 $D=0
M76 vss 153 150 vss n12ll L=6e-08 W=7e-07 $X=6815 $Y=11400 $D=0
M77 vss 148 155 vss n12ll L=6e-08 W=5e-07 $X=6925 $Y=2575 $D=0
M78 151 121 149 vss n12ll L=6e-08 W=2.5e-06 $X=6945 $Y=17190 $D=0
M79 153 A[7] 362 vss n12ll L=6e-08 W=4e-07 $X=6970 $Y=7215 $D=0
M80 151 152 363 vss n12ll L=6e-08 W=1.495e-06 $X=6970 $Y=12950 $D=0
M81 vss 149 PXA[1] vss n12ll L=6e-08 W=1.5e-06 $X=7090 $Y=24740 $D=0
M82 154 150 vss vss n12ll L=6e-08 W=7e-07 $X=7105 $Y=11400 $D=0
M83 155 148 vss vss n12ll L=6e-08 W=5e-07 $X=7215 $Y=2575 $D=0
M84 155 121 163 vss n12ll L=6e-08 W=1.25e-06 $X=7875 $Y=2555 $D=0
M85 163 121 155 vss n12ll L=6e-08 W=1.25e-06 $X=8165 $Y=2555 $D=0
M86 160 158 vss vss n12ll L=6e-08 W=4e-07 $X=8685 $Y=25185 $D=0
M87 FCKX[3] 160 180 vss n12ll L=6e-08 W=1.25e-06 $X=8685 $Y=29105 $D=0
M88 vss vss A[5] vss n12ll L=6e-08 W=2e-07 $X=8740 $Y=14765 $D=0
M89 161 121 158 vss n12ll L=6e-08 W=5e-07 $X=8845 $Y=21145 $D=0
M90 vss 160 158 vss n12ll L=6e-07 W=1.2e-07 $X=8935 $Y=26510 $D=0
M91 vss 158 160 vss n12ll L=6e-08 W=4e-07 $X=8975 $Y=25185 $D=0
M92 180 160 FCKX[3] vss n12ll L=6e-08 W=1.25e-06 $X=8975 $Y=29105 $D=0
M93 A[3] vss vss vss n12ll L=6e-08 W=2e-07 $X=9050 $Y=14765 $D=0
M94 364 159 161 vss n12ll L=6e-08 W=1e-06 $X=9075 $Y=19570 $D=0
M95 158 121 161 vss n12ll L=6e-08 W=5e-07 $X=9115 $Y=21145 $D=0
M96 160 158 vss vss n12ll L=6e-08 W=4e-07 $X=9265 $Y=25185 $D=0
M97 FCKX[3] 160 180 vss n12ll L=6e-08 W=1.25e-06 $X=9265 $Y=29105 $D=0
M98 365 162 364 vss n12ll L=6e-08 W=1e-06 $X=9315 $Y=19570 $D=0
M99 161 121 158 vss n12ll L=6e-08 W=5e-07 $X=9395 $Y=21145 $D=0
M100 174 199 vss vss n12ll L=6e-08 W=5e-07 $X=9465 $Y=15160 $D=0
M101 vss 174 365 vss n12ll L=6e-08 W=1e-06 $X=9555 $Y=19570 $D=0
M102 vss 158 160 vss n12ll L=6e-08 W=4e-07 $X=9555 $Y=25185 $D=0
M103 180 160 FCKX[3] vss n12ll L=6e-08 W=1.25e-06 $X=9555 $Y=29105 $D=0
M104 vss 199 174 vss n12ll L=6e-08 W=5e-07 $X=9755 $Y=15160 $D=0
M105 vss ZASX 163 vss n12ll L=6e-07 W=1.2e-07 $X=9795 $Y=2975 $D=0
M106 ZASX 163 vss vss n12ll L=6e-08 W=2.5e-06 $X=9815 $Y=5535 $D=0
M107 366 174 vss vss n12ll L=6e-08 W=1e-06 $X=9845 $Y=19570 $D=0
M108 164 166 vss vss n12ll L=6e-08 W=4e-07 $X=9845 $Y=25185 $D=0
M109 FCKX[2] 164 180 vss n12ll L=6e-08 W=1.25e-06 $X=9845 $Y=29105 $D=0
M110 166 164 vss vss n12ll L=6e-07 W=1.2e-07 $X=9925 $Y=26510 $D=0
M111 166 121 165 vss n12ll L=6e-08 W=5e-07 $X=10005 $Y=21145 $D=0
M112 199 168 vss vss n12ll L=6e-08 W=5e-07 $X=10045 $Y=15160 $D=0
M113 367 162 366 vss n12ll L=6e-08 W=1e-06 $X=10085 $Y=19570 $D=0
M114 vss 163 ZASX vss n12ll L=6e-08 W=2.5e-06 $X=10105 $Y=5535 $D=0
M115 vss 166 164 vss n12ll L=6e-08 W=4e-07 $X=10135 $Y=25185 $D=0
M116 180 164 FCKX[2] vss n12ll L=6e-08 W=1.25e-06 $X=10135 $Y=29105 $D=0
M117 165 121 166 vss n12ll L=6e-08 W=5e-07 $X=10285 $Y=21145 $D=0
M118 165 167 367 vss n12ll L=6e-08 W=1e-06 $X=10325 $Y=19570 $D=0
M119 vss 168 199 vss n12ll L=6e-08 W=5e-07 $X=10335 $Y=15160 $D=0
M120 ZAS 170 vss vss n12ll L=6e-08 W=2.5e-06 $X=10395 $Y=5535 $D=0
M121 164 166 vss vss n12ll L=6e-08 W=4e-07 $X=10425 $Y=25185 $D=0
M122 FCKX[2] 164 180 vss n12ll L=6e-08 W=1.25e-06 $X=10425 $Y=29105 $D=0
M123 166 121 165 vss n12ll L=6e-08 W=5e-07 $X=10555 $Y=21145 $D=0
M124 vss 170 ZAS vss n12ll L=6e-08 W=2.5e-06 $X=10685 $Y=5535 $D=0
M125 vss 166 164 vss n12ll L=6e-08 W=4e-07 $X=10715 $Y=25185 $D=0
M126 180 164 FCKX[2] vss n12ll L=6e-08 W=1.25e-06 $X=10715 $Y=29105 $D=0
M127 368 A[5] 168 vss n12ll L=6e-08 W=4e-07 $X=10965 $Y=15160 $D=0
M128 vss vss CLK vss n12ll L=6e-08 W=2e-07 $X=10985 $Y=4535 $D=0
M129 172 169 vss vss n12ll L=6e-08 W=4e-07 $X=11005 $Y=25185 $D=0
M130 FCKX[0] 172 180 vss n12ll L=6e-08 W=1.25e-06 $X=11005 $Y=29105 $D=0
M131 170 163 vss vss n12ll L=6e-08 W=1e-06 $X=11035 $Y=7035 $D=0
M132 171 CLK vss vss n12ll L=6e-08 W=4e-07 $X=11055 $Y=2915 $D=0
M133 173 121 169 vss n12ll L=6e-08 W=5e-07 $X=11165 $Y=21145 $D=0
M134 vss vdd 368 vss n12ll L=3e-07 W=4e-07 $X=11245 $Y=15160 $D=0
M135 vss 172 169 vss n12ll L=6e-07 W=1.2e-07 $X=11255 $Y=26510 $D=0
M136 vss 169 172 vss n12ll L=6e-08 W=4e-07 $X=11295 $Y=25185 $D=0
M137 180 172 FCKX[0] vss n12ll L=6e-08 W=1.25e-06 $X=11295 $Y=29105 $D=0
M138 369 167 173 vss n12ll L=6e-08 W=1e-06 $X=11395 $Y=19570 $D=0
M139 169 121 173 vss n12ll L=6e-08 W=5e-07 $X=11435 $Y=21145 $D=0
M140 172 169 vss vss n12ll L=6e-08 W=4e-07 $X=11585 $Y=25185 $D=0
M141 FCKX[0] 172 180 vss n12ll L=6e-08 W=1.25e-06 $X=11585 $Y=29105 $D=0
M142 370 207 369 vss n12ll L=6e-08 W=1e-06 $X=11635 $Y=19570 $D=0
M143 173 121 169 vss n12ll L=6e-08 W=5e-07 $X=11715 $Y=21145 $D=0
M144 vss vss CEN vss n12ll L=6e-08 W=2e-07 $X=11735 $Y=2910 $D=0
M145 vss 174 370 vss n12ll L=6e-08 W=1e-06 $X=11875 $Y=19570 $D=0
M146 vss 169 172 vss n12ll L=6e-08 W=4e-07 $X=11875 $Y=25185 $D=0
M147 180 172 FCKX[0] vss n12ll L=6e-08 W=1.25e-06 $X=11875 $Y=29105 $D=0
M148 vss vss vss vss n12ll L=1e-06 W=1e-06 $X=11940 $Y=4720 $D=0
M149 vss vss vss vss n12ll L=1e-06 W=1e-06 $X=11940 $Y=6030 $D=0
M150 371 171 vss vss n12ll L=6e-08 W=1e-06 $X=12075 $Y=2910 $D=0
M151 372 174 vss vss n12ll L=6e-08 W=1e-06 $X=12165 $Y=19570 $D=0
M152 176 177 vss vss n12ll L=6e-08 W=4e-07 $X=12165 $Y=25185 $D=0
M153 FCKX[1] 176 180 vss n12ll L=6e-08 W=1.25e-06 $X=12165 $Y=29105 $D=0
M154 177 176 vss vss n12ll L=6e-07 W=1.2e-07 $X=12245 $Y=26510 $D=0
M155 175 CEN 371 vss n12ll L=6e-08 W=1e-06 $X=12295 $Y=2910 $D=0
M156 177 121 178 vss n12ll L=6e-08 W=5e-07 $X=12325 $Y=21145 $D=0
M157 181 179 vss vss n12ll L=6e-08 W=1.25e-06 $X=12330 $Y=13140 $D=0
M158 373 207 372 vss n12ll L=6e-08 W=1e-06 $X=12405 $Y=19570 $D=0
M159 vss 177 176 vss n12ll L=6e-08 W=4e-07 $X=12455 $Y=25185 $D=0
M160 180 176 FCKX[1] vss n12ll L=6e-08 W=1.25e-06 $X=12455 $Y=29105 $D=0
M161 178 121 177 vss n12ll L=6e-08 W=5e-07 $X=12605 $Y=21145 $D=0
M162 374 vdd vss vss n12ll L=3e-07 W=4e-07 $X=12615 $Y=15160 $D=0
M163 vss 179 181 vss n12ll L=6e-08 W=1.25e-06 $X=12620 $Y=13140 $D=0
M164 178 159 373 vss n12ll L=6e-08 W=1e-06 $X=12645 $Y=19570 $D=0
M165 176 177 vss vss n12ll L=6e-08 W=4e-07 $X=12745 $Y=25185 $D=0
M166 FCKX[1] 176 180 vss n12ll L=6e-08 W=1.25e-06 $X=12745 $Y=29105 $D=0
M167 vss 184 175 vss n12ll L=6e-07 W=1.2e-07 $X=12810 $Y=3200 $D=0
M168 177 121 178 vss n12ll L=6e-08 W=5e-07 $X=12875 $Y=21145 $D=0
M169 179 DBL vss vss n12ll L=6e-08 W=8e-07 $X=12910 $Y=13140 $D=0
M170 vss 177 176 vss n12ll L=6e-08 W=4e-07 $X=13035 $Y=25185 $D=0
M171 180 176 FCKX[1] vss n12ll L=6e-08 W=1.25e-06 $X=13035 $Y=29105 $D=0
M172 183 A[3] 374 vss n12ll L=6e-08 W=4e-07 $X=13135 $Y=15160 $D=0
M173 185 182 vss vss n12ll L=6e-08 W=4e-07 $X=13325 $Y=25185 $D=0
M174 FCKX[7] 185 180 vss n12ll L=6e-08 W=1.25e-06 $X=13325 $Y=29105 $D=0
M175 186 121 182 vss n12ll L=6e-08 W=5e-07 $X=13485 $Y=21145 $D=0
M176 vss 175 184 vss n12ll L=6e-08 W=4e-07 $X=13560 $Y=2910 $D=0
M177 vss 185 182 vss n12ll L=6e-07 W=1.2e-07 $X=13575 $Y=26510 $D=0
M178 vss 182 185 vss n12ll L=6e-08 W=4e-07 $X=13615 $Y=25185 $D=0
M179 180 185 FCKX[7] vss n12ll L=6e-08 W=1.25e-06 $X=13615 $Y=29105 $D=0
M180 205 CLK 202 vss n12ll L=6e-08 W=4e-06 $X=13620 $Y=4340 $D=0
M181 EMCLK 187 vss vss n12ll L=6e-08 W=6.05e-07 $X=13690 $Y=13230 $D=0
M182 375 159 186 vss n12ll L=6e-08 W=1e-06 $X=13715 $Y=19570 $D=0
M183 182 121 186 vss n12ll L=6e-08 W=5e-07 $X=13755 $Y=21145 $D=0
M184 159 183 vss vss n12ll L=6e-08 W=5e-07 $X=13765 $Y=15160 $D=0
M185 188 184 vss vss n12ll L=6e-08 W=5e-07 $X=13850 $Y=2910 $D=0
M186 185 182 vss vss n12ll L=6e-08 W=4e-07 $X=13905 $Y=25185 $D=0
M187 FCKX[7] 185 180 vss n12ll L=6e-08 W=1.25e-06 $X=13905 $Y=29105 $D=0
M188 202 CLK 205 vss n12ll L=6e-08 W=4e-06 $X=13910 $Y=4340 $D=0
M189 376 162 375 vss n12ll L=6e-08 W=1e-06 $X=13955 $Y=19570 $D=0
M190 vss 187 EMCLK vss n12ll L=6e-08 W=6.05e-07 $X=13980 $Y=13230 $D=0
M191 186 121 182 vss n12ll L=6e-08 W=5e-07 $X=14035 $Y=21145 $D=0
M192 vss 183 159 vss n12ll L=6e-08 W=5e-07 $X=14055 $Y=15160 $D=0
M193 vss CLK 188 vss n12ll L=6e-08 W=5e-07 $X=14140 $Y=2910 $D=0
M194 vss 199 376 vss n12ll L=6e-08 W=1e-06 $X=14195 $Y=19570 $D=0
M195 vss 182 185 vss n12ll L=6e-08 W=4e-07 $X=14195 $Y=25185 $D=0
M196 180 185 FCKX[7] vss n12ll L=6e-08 W=1.25e-06 $X=14195 $Y=29105 $D=0
M197 205 CLK 202 vss n12ll L=6e-08 W=4e-06 $X=14200 $Y=4340 $D=0
M198 167 159 vss vss n12ll L=6e-08 W=5e-07 $X=14345 $Y=15160 $D=0
M199 180 129 216 vss n12ll L=6e-08 W=1e-06 $X=14475 $Y=33415 $D=0
M200 217 129 180 vss n12ll L=6e-08 W=1e-06 $X=14475 $Y=33685 $D=0
M201 377 199 vss vss n12ll L=6e-08 W=1e-06 $X=14485 $Y=19570 $D=0
M202 189 191 vss vss n12ll L=6e-08 W=4e-07 $X=14485 $Y=25185 $D=0
M203 FCKX[6] 189 180 vss n12ll L=6e-08 W=1.25e-06 $X=14485 $Y=29105 $D=0
M204 202 CLK 205 vss n12ll L=6e-08 W=4e-06 $X=14490 $Y=4340 $D=0
M205 191 189 vss vss n12ll L=6e-07 W=1.2e-07 $X=14565 $Y=26510 $D=0
M206 vss 159 167 vss n12ll L=6e-08 W=5e-07 $X=14635 $Y=15160 $D=0
M207 191 121 190 vss n12ll L=6e-08 W=5e-07 $X=14645 $Y=21145 $D=0
M208 378 162 377 vss n12ll L=6e-08 W=1e-06 $X=14725 $Y=19570 $D=0
M209 vss 192 187 vss n12ll L=6e-08 W=4e-07 $X=14745 $Y=13245 $D=0
M210 vss 191 189 vss n12ll L=6e-08 W=4e-07 $X=14775 $Y=25185 $D=0
M211 180 189 FCKX[6] vss n12ll L=6e-08 W=1.25e-06 $X=14775 $Y=29105 $D=0
M212 205 CLK 202 vss n12ll L=6e-08 W=4e-06 $X=14780 $Y=4340 $D=0
M213 vss 188 193 vss n12ll L=6e-08 W=5e-07 $X=14830 $Y=2835 $D=0
M214 190 121 191 vss n12ll L=6e-08 W=5e-07 $X=14925 $Y=21145 $D=0
M215 190 167 378 vss n12ll L=6e-08 W=1e-06 $X=14965 $Y=19570 $D=0
M216 192 197 vss vss n12ll L=6e-08 W=4e-07 $X=15035 $Y=13245 $D=0
M217 189 191 vss vss n12ll L=6e-08 W=4e-07 $X=15065 $Y=25185 $D=0
M218 FCKX[6] 189 180 vss n12ll L=6e-08 W=1.25e-06 $X=15065 $Y=29105 $D=0
M219 194 193 vss vss n12ll L=6e-08 W=7.5e-07 $X=15180 $Y=2835 $D=0
M220 191 121 190 vss n12ll L=6e-08 W=5e-07 $X=15195 $Y=21145 $D=0
M221 vss 191 189 vss n12ll L=6e-08 W=4e-07 $X=15355 $Y=25185 $D=0
M222 180 189 FCKX[6] vss n12ll L=6e-08 W=1.25e-06 $X=15355 $Y=29105 $D=0
M223 205 194 vss vss n12ll L=6e-08 W=2.5e-06 $X=15440 $Y=5495 $D=0
M224 vss 193 194 vss n12ll L=6e-08 W=7.5e-07 $X=15470 $Y=2835 $D=0
M225 379 vdd vss vss n12ll L=3e-07 W=4e-07 $X=15515 $Y=15160 $D=0
M226 196 195 vss vss n12ll L=6e-08 W=4e-07 $X=15645 $Y=25185 $D=0
M227 FCKX[4] 196 180 vss n12ll L=6e-08 W=1.25e-06 $X=15645 $Y=29105 $D=0
M228 vss 194 205 vss n12ll L=6e-08 W=2.5e-06 $X=15730 $Y=5495 $D=0
M229 198 121 195 vss n12ll L=6e-08 W=5e-07 $X=15805 $Y=21145 $D=0
M230 221 215 vss vss n12ll L=6e-08 W=1.5e-06 $X=15870 $Y=2835 $D=0
M231 vss 196 195 vss n12ll L=6e-07 W=1.2e-07 $X=15895 $Y=26510 $D=0
M232 vss 195 196 vss n12ll L=6e-08 W=4e-07 $X=15935 $Y=25185 $D=0
M233 180 196 FCKX[4] vss n12ll L=6e-08 W=1.25e-06 $X=15935 $Y=29105 $D=0
M234 205 194 vss vss n12ll L=6e-08 W=2.5e-06 $X=16020 $Y=5495 $D=0
M235 200 A[4] 379 vss n12ll L=6e-08 W=4e-07 $X=16035 $Y=15160 $D=0
M236 380 167 198 vss n12ll L=6e-08 W=1e-06 $X=16035 $Y=19570 $D=0
M237 195 121 198 vss n12ll L=6e-08 W=5e-07 $X=16075 $Y=21145 $D=0
M238 vss 215 221 vss n12ll L=6e-08 W=1.5e-06 $X=16185 $Y=2835 $D=0
M239 196 195 vss vss n12ll L=6e-08 W=4e-07 $X=16225 $Y=25185 $D=0
M240 FCKX[4] 196 180 vss n12ll L=6e-08 W=1.25e-06 $X=16225 $Y=29105 $D=0
M241 381 207 380 vss n12ll L=6e-08 W=1e-06 $X=16275 $Y=19570 $D=0
M242 vss 194 205 vss n12ll L=6e-08 W=2.5e-06 $X=16310 $Y=5495 $D=0
M243 vss 201 197 vss n12ll L=6e-08 W=4e-07 $X=16320 $Y=13245 $D=0
M244 198 121 195 vss n12ll L=6e-08 W=5e-07 $X=16355 $Y=21145 $D=0
M245 vss 199 381 vss n12ll L=6e-08 W=1e-06 $X=16515 $Y=19570 $D=0
M246 vss 195 196 vss n12ll L=6e-08 W=4e-07 $X=16515 $Y=25185 $D=0
M247 180 196 FCKX[4] vss n12ll L=6e-08 W=1.25e-06 $X=16515 $Y=29105 $D=0
M248 204 251 vss vss n12ll L=6e-08 W=7.5e-07 $X=16540 $Y=2835 $D=0
M249 205 194 vss vss n12ll L=6e-08 W=2.5e-06 $X=16600 $Y=5495 $D=0
M250 162 200 vss vss n12ll L=6e-08 W=5e-07 $X=16665 $Y=15160 $D=0
M251 201 202 vss vss n12ll L=6e-08 W=7e-07 $X=16670 $Y=13245 $D=0
M252 382 199 vss vss n12ll L=6e-08 W=1e-06 $X=16805 $Y=19570 $D=0
M253 206 208 vss vss n12ll L=6e-08 W=4e-07 $X=16805 $Y=25185 $D=0
M254 FCKX[5] 206 180 vss n12ll L=6e-08 W=1.25e-06 $X=16805 $Y=29105 $D=0
M255 vss 211 204 vss n12ll L=6e-08 W=7.5e-07 $X=16830 $Y=2835 $D=0
M256 208 206 vss vss n12ll L=6e-07 W=1.2e-07 $X=16885 $Y=26510 $D=0
M257 vss 194 205 vss n12ll L=6e-08 W=2.5e-06 $X=16890 $Y=5495 $D=0
M258 vss 200 162 vss n12ll L=6e-08 W=5e-07 $X=16955 $Y=15160 $D=0
M259 208 121 210 vss n12ll L=6e-08 W=5e-07 $X=16965 $Y=21145 $D=0
M260 383 207 382 vss n12ll L=6e-08 W=1e-06 $X=17045 $Y=19570 $D=0
M261 vss 208 206 vss n12ll L=6e-08 W=4e-07 $X=17095 $Y=25185 $D=0
M262 180 206 FCKX[5] vss n12ll L=6e-08 W=1.25e-06 $X=17095 $Y=29105 $D=0
M263 204 211 vss vss n12ll L=6e-08 W=7.5e-07 $X=17120 $Y=2835 $D=0
M264 205 194 vss vss n12ll L=6e-08 W=2.5e-06 $X=17180 $Y=5495 $D=0
M265 207 162 vss vss n12ll L=6e-08 W=5e-07 $X=17245 $Y=15160 $D=0
M266 210 121 208 vss n12ll L=6e-08 W=5e-07 $X=17245 $Y=21145 $D=0
M267 210 159 383 vss n12ll L=6e-08 W=1e-06 $X=17285 $Y=19570 $D=0
M268 206 208 vss vss n12ll L=6e-08 W=4e-07 $X=17385 $Y=25185 $D=0
M269 FCKX[5] 206 180 vss n12ll L=6e-08 W=1.25e-06 $X=17385 $Y=29105 $D=0
M270 vss 251 204 vss n12ll L=6e-08 W=7.5e-07 $X=17410 $Y=2835 $D=0
M271 vss 194 205 vss n12ll L=6e-08 W=2.5e-06 $X=17470 $Y=5495 $D=0
M272 208 121 210 vss n12ll L=6e-08 W=5e-07 $X=17515 $Y=21145 $D=0
M273 vss 162 207 vss n12ll L=6e-08 W=5e-07 $X=17535 $Y=15160 $D=0
M274 vss 208 206 vss n12ll L=6e-08 W=4e-07 $X=17675 $Y=25185 $D=0
M275 180 206 FCKX[5] vss n12ll L=6e-08 W=1.25e-06 $X=17675 $Y=29105 $D=0
M276 215 209 vss vss n12ll L=6e-08 W=2.5e-06 $X=17760 $Y=5495 $D=0
M277 vss vss A[4] vss n12ll L=6e-08 W=2e-07 $X=17940 $Y=14820 $D=0
M278 214 212 vss vss n12ll L=6e-08 W=4e-07 $X=17965 $Y=25185 $D=0
M279 YX[3] 214 180 vss n12ll L=6e-08 W=1.25e-06 $X=17965 $Y=29105 $D=0
M280 vss 251 215 vss n12ll L=6e-08 W=2.5e-06 $X=18050 $Y=5495 $D=0
M281 vss 219 211 vss n12ll L=2e-07 W=4e-07 $X=18100 $Y=2860 $D=0
M282 218 121 212 vss n12ll L=6e-08 W=5e-07 $X=18125 $Y=21145 $D=0
M283 vss 214 212 vss n12ll L=6e-07 W=1.2e-07 $X=18215 $Y=26510 $D=0
M284 A[2] vss vss vss n12ll L=6e-08 W=2e-07 $X=18250 $Y=14820 $D=0
M285 vss 212 214 vss n12ll L=6e-08 W=4e-07 $X=18255 $Y=25185 $D=0
M286 180 214 YX[3] vss n12ll L=6e-08 W=1.25e-06 $X=18255 $Y=29105 $D=0
M287 120 215 vss vss n12ll L=6e-08 W=2.5e-06 $X=18340 $Y=5495 $D=0
M288 384 213 218 vss n12ll L=6e-08 W=1e-06 $X=18355 $Y=19570 $D=0
M289 212 121 218 vss n12ll L=6e-08 W=5e-07 $X=18395 $Y=21145 $D=0
M290 214 212 vss vss n12ll L=6e-08 W=4e-07 $X=18545 $Y=25185 $D=0
M291 YX[3] 214 180 vss n12ll L=6e-08 W=1.25e-06 $X=18545 $Y=29105 $D=0
M292 219 251 vss vss n12ll L=2e-07 W=4e-07 $X=18590 $Y=2860 $D=0
M293 385 220 384 vss n12ll L=6e-08 W=1e-06 $X=18595 $Y=19570 $D=0
M294 vss 215 120 vss n12ll L=6e-08 W=2.5e-06 $X=18630 $Y=5495 $D=0
M295 218 121 212 vss n12ll L=6e-08 W=5e-07 $X=18675 $Y=21145 $D=0
M296 231 249 vss vss n12ll L=6e-08 W=5e-07 $X=18745 $Y=15160 $D=0
M297 vss 216 RWLL vss n12ll L=6e-08 W=2e-06 $X=18775 $Y=33415 $D=0
M298 RWLR 217 vss vss n12ll L=6e-08 W=2e-06 $X=18775 $Y=33685 $D=0
M299 vss 231 385 vss n12ll L=6e-08 W=1e-06 $X=18835 $Y=19570 $D=0
M300 vss 212 214 vss n12ll L=6e-08 W=4e-07 $X=18835 $Y=25185 $D=0
M301 180 214 YX[3] vss n12ll L=6e-08 W=1.25e-06 $X=18835 $Y=29105 $D=0
M302 DCTRCLK 215 vss vss n12ll L=6e-08 W=2.5e-06 $X=18920 $Y=5495 $D=0
M303 vss 249 231 vss n12ll L=6e-08 W=5e-07 $X=19035 $Y=15160 $D=0
M304 386 231 vss vss n12ll L=6e-08 W=1e-06 $X=19125 $Y=19570 $D=0
M305 222 224 vss vss n12ll L=6e-08 W=4e-07 $X=19125 $Y=25185 $D=0
M306 YX[2] 222 180 vss n12ll L=6e-08 W=1.25e-06 $X=19125 $Y=29105 $D=0
M307 224 222 vss vss n12ll L=6e-07 W=1.2e-07 $X=19205 $Y=26510 $D=0
M308 vss 215 DCTRCLK vss n12ll L=6e-08 W=2.5e-06 $X=19210 $Y=5495 $D=0
M309 224 121 223 vss n12ll L=6e-08 W=5e-07 $X=19285 $Y=21145 $D=0
M310 249 226 vss vss n12ll L=6e-08 W=5e-07 $X=19325 $Y=15160 $D=0
M311 387 220 386 vss n12ll L=6e-08 W=1e-06 $X=19365 $Y=19570 $D=0
M312 vss 228 209 vss n12ll L=2e-07 W=4e-07 $X=19410 $Y=2745 $D=0
M313 vss 224 222 vss n12ll L=6e-08 W=4e-07 $X=19415 $Y=25185 $D=0
M314 180 222 YX[2] vss n12ll L=6e-08 W=1.25e-06 $X=19415 $Y=29105 $D=0
M315 121 120 vss vss n12ll L=6e-08 W=2.5e-06 $X=19500 $Y=5495 $D=0
M316 223 121 224 vss n12ll L=6e-08 W=5e-07 $X=19565 $Y=21145 $D=0
M317 223 225 387 vss n12ll L=6e-08 W=1e-06 $X=19605 $Y=19570 $D=0
M318 vss 226 249 vss n12ll L=6e-08 W=5e-07 $X=19615 $Y=15160 $D=0
M319 222 224 vss vss n12ll L=6e-08 W=4e-07 $X=19705 $Y=25185 $D=0
M320 YX[2] 222 180 vss n12ll L=6e-08 W=1.25e-06 $X=19705 $Y=29105 $D=0
M321 vss 120 121 vss n12ll L=6e-08 W=2.5e-06 $X=19790 $Y=5495 $D=0
M322 224 121 223 vss n12ll L=6e-08 W=5e-07 $X=19835 $Y=21145 $D=0
M323 228 vss vss vss n12ll L=2e-07 W=4e-07 $X=19900 $Y=2745 $D=0
M324 vss 224 222 vss n12ll L=6e-08 W=4e-07 $X=19995 $Y=25185 $D=0
M325 180 222 YX[2] vss n12ll L=6e-08 W=1.25e-06 $X=19995 $Y=29105 $D=0
M326 vss 251 202 vss n12ll L=1e-06 W=1.2e-07 $X=20075 $Y=3695 $D=0
M327 DCTRCLKX 221 vss vss n12ll L=6e-08 W=2.5e-06 $X=20080 $Y=5495 $D=0
M328 388 A[2] 226 vss n12ll L=6e-08 W=4e-07 $X=20245 $Y=15160 $D=0
M329 229 227 vss vss n12ll L=6e-08 W=4e-07 $X=20285 $Y=25185 $D=0
M330 YX[0] 229 180 vss n12ll L=6e-08 W=1.25e-06 $X=20285 $Y=29105 $D=0
M331 vss vss WEN vss n12ll L=6e-08 W=2e-07 $X=20360 $Y=4745 $D=0
M332 vss 221 DCTRCLKX vss n12ll L=6e-08 W=2.5e-06 $X=20370 $Y=5495 $D=0
M333 vss 251 228 vss n12ll L=2e-07 W=4e-07 $X=20390 $Y=2745 $D=0
M334 230 121 227 vss n12ll L=6e-08 W=5e-07 $X=20445 $Y=21145 $D=0
M335 vss vdd 388 vss n12ll L=3e-07 W=4e-07 $X=20525 $Y=15160 $D=0
M336 vss 229 227 vss n12ll L=6e-07 W=1.2e-07 $X=20535 $Y=26510 $D=0
M337 vss 227 229 vss n12ll L=6e-08 W=4e-07 $X=20575 $Y=25185 $D=0
M338 180 229 YX[0] vss n12ll L=6e-08 W=1.25e-06 $X=20575 $Y=29105 $D=0
M339 SACK4 204 vss vss n12ll L=6e-08 W=2.5e-06 $X=20660 $Y=5495 $D=0
M340 389 225 230 vss n12ll L=6e-08 W=1e-06 $X=20675 $Y=19570 $D=0
M341 227 121 230 vss n12ll L=6e-08 W=5e-07 $X=20715 $Y=21145 $D=0
M342 229 227 vss vss n12ll L=6e-08 W=4e-07 $X=20865 $Y=25185 $D=0
M343 YX[0] 229 180 vss n12ll L=6e-08 W=1.25e-06 $X=20865 $Y=29105 $D=0
M344 390 254 389 vss n12ll L=6e-08 W=1e-06 $X=20915 $Y=19570 $D=0
M345 vss 204 SACK4 vss n12ll L=6e-08 W=2.5e-06 $X=20950 $Y=5495 $D=0
M346 230 121 227 vss n12ll L=6e-08 W=5e-07 $X=20995 $Y=21145 $D=0
M347 vss 231 390 vss n12ll L=6e-08 W=1e-06 $X=21155 $Y=19570 $D=0
M348 vss 227 229 vss n12ll L=6e-08 W=4e-07 $X=21155 $Y=25185 $D=0
M349 180 229 YX[0] vss n12ll L=6e-08 W=1.25e-06 $X=21155 $Y=29105 $D=0
M350 vss WEN 232 vss n12ll L=6e-08 W=4e-07 $X=21180 $Y=2745 $D=0
M351 251 202 vss vss n12ll L=6e-08 W=2.5e-06 $X=21240 $Y=5495 $D=0
M352 391 231 vss vss n12ll L=6e-08 W=1e-06 $X=21445 $Y=19570 $D=0
M353 233 234 vss vss n12ll L=6e-08 W=4e-07 $X=21445 $Y=25185 $D=0
M354 YX[1] 233 180 vss n12ll L=6e-08 W=1.25e-06 $X=21445 $Y=29105 $D=0
M355 236 232 vss vss n12ll L=3e-07 W=4e-07 $X=21500 $Y=2745 $D=0
M356 234 233 vss vss n12ll L=6e-07 W=1.2e-07 $X=21525 $Y=26510 $D=0
M357 vss 202 251 vss n12ll L=6e-08 W=2.5e-06 $X=21530 $Y=5495 $D=0
M358 234 121 235 vss n12ll L=6e-08 W=5e-07 $X=21605 $Y=21145 $D=0
M359 392 254 391 vss n12ll L=6e-08 W=1e-06 $X=21685 $Y=19570 $D=0
M360 vss 234 233 vss n12ll L=6e-08 W=4e-07 $X=21735 $Y=25185 $D=0
M361 180 233 YX[1] vss n12ll L=6e-08 W=1.25e-06 $X=21735 $Y=29105 $D=0
M362 251 202 vss vss n12ll L=6e-08 W=2.5e-06 $X=21820 $Y=5495 $D=0
M363 235 121 234 vss n12ll L=6e-08 W=5e-07 $X=21885 $Y=21145 $D=0
M364 393 vdd vss vss n12ll L=3e-07 W=4e-07 $X=21895 $Y=15160 $D=0
M365 235 213 392 vss n12ll L=6e-08 W=1e-06 $X=21925 $Y=19570 $D=0
M366 233 234 vss vss n12ll L=6e-08 W=4e-07 $X=22025 $Y=25185 $D=0
M367 YX[1] 233 180 vss n12ll L=6e-08 W=1.25e-06 $X=22025 $Y=29105 $D=0
M368 vss 202 251 vss n12ll L=6e-08 W=2.5e-06 $X=22110 $Y=5495 $D=0
M369 234 121 235 vss n12ll L=6e-08 W=5e-07 $X=22155 $Y=21145 $D=0
M370 vss 234 233 vss n12ll L=6e-08 W=4e-07 $X=22315 $Y=25185 $D=0
M371 180 233 YX[1] vss n12ll L=6e-08 W=1.25e-06 $X=22315 $Y=29105 $D=0
M372 SACK1 251 vss vss n12ll L=6e-08 W=2.5e-06 $X=22400 $Y=5495 $D=0
M373 238 A[0] 393 vss n12ll L=6e-08 W=4e-07 $X=22415 $Y=15160 $D=0
M374 vss 236 239 vss n12ll L=2e-07 W=4e-07 $X=22460 $Y=2795 $D=0
M375 241 237 vss vss n12ll L=6e-08 W=4e-07 $X=22605 $Y=25185 $D=0
M376 YX[7] 241 180 vss n12ll L=6e-08 W=1.25e-06 $X=22605 $Y=29105 $D=0
M377 vss 251 SACK1 vss n12ll L=6e-08 W=2.5e-06 $X=22690 $Y=5495 $D=0
M378 242 121 237 vss n12ll L=6e-08 W=5e-07 $X=22765 $Y=21145 $D=0
M379 vss 241 237 vss n12ll L=6e-07 W=1.2e-07 $X=22855 $Y=26510 $D=0
M380 vss 237 241 vss n12ll L=6e-08 W=4e-07 $X=22895 $Y=25185 $D=0
M381 180 241 YX[7] vss n12ll L=6e-08 W=1.25e-06 $X=22895 $Y=29105 $D=0
M382 180 251 vss vss n12ll L=6e-08 W=2.5e-06 $X=22980 $Y=5495 $D=0
M383 240 239 vss vss n12ll L=6e-08 W=1e-06 $X=22995 $Y=2795 $D=0
M384 394 213 242 vss n12ll L=6e-08 W=1e-06 $X=22995 $Y=19570 $D=0
M385 237 121 242 vss n12ll L=6e-08 W=5e-07 $X=23035 $Y=21145 $D=0
M386 213 238 vss vss n12ll L=6e-08 W=5e-07 $X=23045 $Y=15160 $D=0
M387 241 237 vss vss n12ll L=6e-08 W=4e-07 $X=23185 $Y=25185 $D=0
M388 YX[7] 241 180 vss n12ll L=6e-08 W=1.25e-06 $X=23185 $Y=29105 $D=0
M389 395 220 394 vss n12ll L=6e-08 W=1e-06 $X=23235 $Y=19570 $D=0
M390 vss 251 180 vss n12ll L=6e-08 W=2.5e-06 $X=23270 $Y=5495 $D=0
M391 257 121 240 vss n12ll L=6e-08 W=1e-06 $X=23285 $Y=2795 $D=0
M392 242 121 237 vss n12ll L=6e-08 W=5e-07 $X=23315 $Y=21145 $D=0
M393 vss 238 213 vss n12ll L=6e-08 W=5e-07 $X=23335 $Y=15160 $D=0
M394 vss 249 395 vss n12ll L=6e-08 W=1e-06 $X=23475 $Y=19570 $D=0
M395 vss 237 241 vss n12ll L=6e-08 W=4e-07 $X=23475 $Y=25185 $D=0
M396 180 241 YX[7] vss n12ll L=6e-08 W=1.25e-06 $X=23475 $Y=29105 $D=0
M397 180 251 vss vss n12ll L=6e-08 W=2.5e-06 $X=23560 $Y=5495 $D=0
M398 225 213 vss vss n12ll L=6e-08 W=5e-07 $X=23625 $Y=15160 $D=0
M399 396 249 vss vss n12ll L=6e-08 W=1e-06 $X=23765 $Y=19570 $D=0
M400 243 245 vss vss n12ll L=6e-08 W=4e-07 $X=23765 $Y=25185 $D=0
M401 YX[6] 243 180 vss n12ll L=6e-08 W=1.25e-06 $X=23765 $Y=29105 $D=0
M402 245 243 vss vss n12ll L=6e-07 W=1.2e-07 $X=23845 $Y=26510 $D=0
M403 vss 251 180 vss n12ll L=6e-08 W=2.5e-06 $X=23850 $Y=5495 $D=0
M404 vss 213 225 vss n12ll L=6e-08 W=5e-07 $X=23915 $Y=15160 $D=0
M405 245 121 244 vss n12ll L=6e-08 W=5e-07 $X=23925 $Y=21145 $D=0
M406 397 220 396 vss n12ll L=6e-08 W=1e-06 $X=24005 $Y=19570 $D=0
M407 vss 245 243 vss n12ll L=6e-08 W=4e-07 $X=24055 $Y=25185 $D=0
M408 180 243 YX[6] vss n12ll L=6e-08 W=1.25e-06 $X=24055 $Y=29105 $D=0
M409 180 251 vss vss n12ll L=6e-08 W=2.5e-06 $X=24140 $Y=5495 $D=0
M410 244 121 245 vss n12ll L=6e-08 W=5e-07 $X=24205 $Y=21145 $D=0
M411 244 225 397 vss n12ll L=6e-08 W=1e-06 $X=24245 $Y=19570 $D=0
M412 243 245 vss vss n12ll L=6e-08 W=4e-07 $X=24345 $Y=25185 $D=0
M413 YX[6] 243 180 vss n12ll L=6e-08 W=1.25e-06 $X=24345 $Y=29105 $D=0
M414 vss vss A[0] vss n12ll L=6e-08 W=2e-07 $X=24395 $Y=14735 $D=0
M415 vss 251 180 vss n12ll L=6e-08 W=2.5e-06 $X=24430 $Y=5495 $D=0
M416 245 121 244 vss n12ll L=6e-08 W=5e-07 $X=24475 $Y=21145 $D=0
M417 vss 245 243 vss n12ll L=6e-08 W=4e-07 $X=24635 $Y=25185 $D=0
M418 180 243 YX[6] vss n12ll L=6e-08 W=1.25e-06 $X=24635 $Y=29105 $D=0
M419 180 251 vss vss n12ll L=6e-08 W=2.5e-06 $X=24720 $Y=5495 $D=0
M420 398 vdd vss vss n12ll L=3e-07 W=4e-07 $X=24795 $Y=15160 $D=0
M421 247 246 vss vss n12ll L=6e-08 W=4e-07 $X=24925 $Y=25185 $D=0
M422 YX[4] 247 180 vss n12ll L=6e-08 W=1.25e-06 $X=24925 $Y=29105 $D=0
M423 vss 251 180 vss n12ll L=6e-08 W=2.5e-06 $X=25010 $Y=5495 $D=0
M424 248 121 246 vss n12ll L=6e-08 W=5e-07 $X=25085 $Y=21145 $D=0
M425 vss 247 246 vss n12ll L=6e-07 W=1.2e-07 $X=25175 $Y=26510 $D=0
M426 vss 246 247 vss n12ll L=6e-08 W=4e-07 $X=25215 $Y=25185 $D=0
M427 180 247 YX[4] vss n12ll L=6e-08 W=1.25e-06 $X=25215 $Y=29105 $D=0
M428 WE 252 vss vss n12ll L=6e-08 W=2.5e-06 $X=25300 $Y=5495 $D=0
M429 250 A[1] 398 vss n12ll L=6e-08 W=4e-07 $X=25315 $Y=15160 $D=0
M430 399 225 248 vss n12ll L=6e-08 W=1e-06 $X=25315 $Y=19570 $D=0
M431 246 121 248 vss n12ll L=6e-08 W=5e-07 $X=25355 $Y=21145 $D=0
M432 247 246 vss vss n12ll L=6e-08 W=4e-07 $X=25505 $Y=25185 $D=0
M433 YX[4] 247 180 vss n12ll L=6e-08 W=1.25e-06 $X=25505 $Y=29105 $D=0
M434 400 254 399 vss n12ll L=6e-08 W=1e-06 $X=25555 $Y=19570 $D=0
M435 vss 252 WE vss n12ll L=6e-08 W=2.5e-06 $X=25590 $Y=5495 $D=0
M436 248 121 246 vss n12ll L=6e-08 W=5e-07 $X=25635 $Y=21145 $D=0
M437 vss vss A[1] vss n12ll L=6e-08 W=2e-07 $X=25725 $Y=14735 $D=0
M438 vss 249 400 vss n12ll L=6e-08 W=1e-06 $X=25795 $Y=19570 $D=0
M439 vss 246 247 vss n12ll L=6e-08 W=4e-07 $X=25795 $Y=25185 $D=0
M440 180 247 YX[4] vss n12ll L=6e-08 W=1.25e-06 $X=25795 $Y=29105 $D=0
M441 401 258 vss vss n12ll L=6e-08 W=3e-06 $X=25880 $Y=4995 $D=0
M442 220 250 vss vss n12ll L=6e-08 W=5e-07 $X=25945 $Y=15160 $D=0
M443 402 249 vss vss n12ll L=6e-08 W=1e-06 $X=26085 $Y=19570 $D=0
M444 253 255 vss vss n12ll L=6e-08 W=4e-07 $X=26085 $Y=25185 $D=0
M445 YX[5] 253 180 vss n12ll L=6e-08 W=1.25e-06 $X=26085 $Y=29105 $D=0
M446 255 253 vss vss n12ll L=6e-07 W=1.2e-07 $X=26165 $Y=26510 $D=0
M447 252 251 401 vss n12ll L=6e-08 W=3e-06 $X=26170 $Y=4995 $D=0
M448 vss 250 220 vss n12ll L=6e-08 W=5e-07 $X=26235 $Y=15160 $D=0
M449 255 121 256 vss n12ll L=6e-08 W=5e-07 $X=26245 $Y=21145 $D=0
M450 403 254 402 vss n12ll L=6e-08 W=1e-06 $X=26325 $Y=19570 $D=0
M451 vss 255 253 vss n12ll L=6e-08 W=4e-07 $X=26375 $Y=25185 $D=0
M452 180 253 YX[5] vss n12ll L=6e-08 W=1.25e-06 $X=26375 $Y=29105 $D=0
M453 254 220 vss vss n12ll L=6e-08 W=5e-07 $X=26525 $Y=15160 $D=0
M454 256 121 255 vss n12ll L=6e-08 W=5e-07 $X=26525 $Y=21145 $D=0
M455 256 213 403 vss n12ll L=6e-08 W=1e-06 $X=26565 $Y=19570 $D=0
M456 253 255 vss vss n12ll L=6e-08 W=4e-07 $X=26665 $Y=25185 $D=0
M457 YX[5] 253 180 vss n12ll L=6e-08 W=1.25e-06 $X=26665 $Y=29105 $D=0
M458 255 121 256 vss n12ll L=6e-08 W=5e-07 $X=26795 $Y=21145 $D=0
M459 vss 220 254 vss n12ll L=6e-08 W=5e-07 $X=26815 $Y=15160 $D=0
M460 vss 257 258 vss n12ll L=6e-08 W=1e-06 $X=26930 $Y=7035 $D=0
M461 vss 255 253 vss n12ll L=6e-08 W=4e-07 $X=26955 $Y=25185 $D=0
M462 180 253 YX[5] vss n12ll L=6e-08 W=1.25e-06 $X=26955 $Y=29105 $D=0
M463 vss 258 257 vss n12ll L=6e-07 W=1.2e-07 $X=26960 $Y=5345 $D=0
M464 410 vss vdd vdd p12ll L=1e-07 W=4e-07 $X=810 $Y=1515 $D=2
M465 99 RDE 410 vdd p12ll L=6e-08 W=4e-07 $X=1110 $Y=1515 $D=2
M466 114 99 vdd vdd p12ll L=6e-08 W=8e-07 $X=1700 $Y=1315 $D=2
M467 124 126 vdd vdd p12ll L=3e-07 W=1.2e-07 $X=1965 $Y=660 $D=2
M468 vdd 114 115 vdd p12ll L=6e-08 W=8e-07 $X=2320 $Y=1315 $D=2
M469 PXB[3] 118 vdd vdd p12ll L=6e-08 W=3.5e-06 $X=2590 $Y=26845 $D=2
M470 119 115 vdd vdd p12ll L=6e-08 W=8e-07 $X=2600 $Y=1315 $D=2
M471 116 135 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=2610 $Y=15140 $D=2
M472 421 A[8] 117 vdd p12ll L=6e-08 W=4e-07 $X=2730 $Y=8445 $D=2
M473 118 120 116 vdd p12ll L=6e-08 W=2.5e-06 $X=2735 $Y=20205 $D=2
M474 123 PXB[2] vdd vdd p12ll L=3e-07 W=1.2e-07 $X=2870 $Y=30975 $D=2
M475 vdd 118 PXB[3] vdd p12ll L=6e-08 W=3.5e-06 $X=2880 $Y=26845 $D=2
M476 vdd 130 116 vdd p12ll L=6e-08 W=1.5e-06 $X=2890 $Y=15140 $D=2
M477 vdd 117 135 vdd p12ll L=6e-08 W=1.4e-06 $X=2925 $Y=9390 $D=2
M478 vdd vdd A[8] vdd p12ll L=6e-08 W=2e-07 $X=2935 $Y=5240 $D=2
M479 vdd vss 421 vdd p12ll L=1e-07 W=4e-07 $X=3045 $Y=8445 $D=2
M480 124 120 119 vdd p12ll L=6e-08 W=1e-06 $X=3060 $Y=1145 $D=2
M481 vdd PXB[3] 118 vdd p12ll L=3e-07 W=1.2e-07 $X=3125 $Y=31630 $D=2
M482 122 130 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=3160 $Y=15140 $D=2
M483 PXB[2] 123 vdd vdd p12ll L=6e-08 W=3.5e-06 $X=3170 $Y=26845 $D=2
M484 125 135 vdd vdd p12ll L=6e-08 W=1.4e-06 $X=3215 $Y=9390 $D=2
M485 122 120 123 vdd p12ll L=6e-08 W=2.5e-06 $X=3315 $Y=20205 $D=2
M486 vdd 125 122 vdd p12ll L=6e-08 W=1.5e-06 $X=3440 $Y=15140 $D=2
M487 vdd 123 PXB[2] vdd p12ll L=6e-08 W=3.5e-06 $X=3460 $Y=26845 $D=2
M488 vdd 124 126 vdd p12ll L=6e-08 W=8e-07 $X=3670 $Y=1315 $D=2
M489 PXB[0] 127 vdd vdd p12ll L=6e-08 W=3.5e-06 $X=3800 $Y=26845 $D=2
M490 128 125 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=3820 $Y=15140 $D=2
M491 132 PXB[1] vdd vdd p12ll L=3e-07 W=1.2e-07 $X=3895 $Y=31630 $D=2
M492 127 120 128 vdd p12ll L=6e-08 W=2.5e-06 $X=3945 $Y=20205 $D=2
M493 129 126 vdd vdd p12ll L=6e-08 W=8e-07 $X=3950 $Y=1315 $D=2
M494 vdd 133 130 vdd p12ll L=6e-08 W=1.4e-06 $X=4045 $Y=9390 $D=2
M495 vdd 127 PXB[0] vdd p12ll L=6e-08 W=3.5e-06 $X=4090 $Y=26845 $D=2
M496 vdd 131 128 vdd p12ll L=6e-08 W=1.5e-06 $X=4100 $Y=15140 $D=2
M497 vdd PXB[0] 127 vdd p12ll L=3e-07 W=1.2e-07 $X=4150 $Y=30975 $D=2
M498 423 vss vdd vdd p12ll L=1e-07 W=4e-07 $X=4195 $Y=8445 $D=2
M499 131 130 vdd vdd p12ll L=6e-08 W=1.4e-06 $X=4335 $Y=9390 $D=2
M500 134 131 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=4370 $Y=15140 $D=2
M501 PXB[1] 132 vdd vdd p12ll L=6e-08 W=3.5e-06 $X=4380 $Y=26845 $D=2
M502 134 120 132 vdd p12ll L=6e-08 W=2.5e-06 $X=4525 $Y=20205 $D=2
M503 133 A[9] 423 vdd p12ll L=6e-08 W=4e-07 $X=4550 $Y=8445 $D=2
M504 vdd 135 134 vdd p12ll L=6e-08 W=1.5e-06 $X=4650 $Y=15140 $D=2
M505 vdd 132 PXB[1] vdd p12ll L=6e-08 W=3.5e-06 $X=4670 $Y=26845 $D=2
M506 vdd vdd A[9] vdd p12ll L=6e-08 W=2e-07 $X=4745 $Y=5260 $D=2
M507 vdd A[6] 137 vdd p12ll L=6e-08 W=4e-07 $X=4975 $Y=1395 $D=2
M508 PXA[3] 139 vdd vdd p12ll L=6e-08 W=3.5e-06 $X=5010 $Y=26845 $D=2
M509 138 152 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=5030 $Y=15140 $D=2
M510 139 120 138 vdd p12ll L=6e-08 W=2.5e-06 $X=5155 $Y=20205 $D=2
M511 424 140 152 vdd p12ll L=6e-08 W=7e-07 $X=5165 $Y=10090 $D=2
M512 142 PXA[2] vdd vdd p12ll L=3e-07 W=1.2e-07 $X=5290 $Y=30975 $D=2
M513 vdd 139 PXA[3] vdd p12ll L=6e-08 W=3.5e-06 $X=5300 $Y=26845 $D=2
M514 vdd 150 138 vdd p12ll L=6e-08 W=1.5e-06 $X=5310 $Y=15140 $D=2
M515 145 137 vdd vdd p12ll L=3e-07 W=4e-07 $X=5335 $Y=1395 $D=2
M516 vdd A[6] 140 vdd p12ll L=6e-08 W=4e-07 $X=5375 $Y=8290 $D=2
M517 vdd RDE 424 vdd p12ll L=6e-08 W=7e-07 $X=5455 $Y=10090 $D=2
M518 vdd PXA[3] 139 vdd p12ll L=3e-07 W=1.2e-07 $X=5545 $Y=31630 $D=2
M519 141 150 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=5580 $Y=15140 $D=2
M520 PXA[2] 142 vdd vdd p12ll L=6e-08 W=3.5e-06 $X=5590 $Y=26845 $D=2
M521 143 140 vdd vdd p12ll L=6e-08 W=4e-07 $X=5655 $Y=8290 $D=2
M522 141 120 142 vdd p12ll L=6e-08 W=2.5e-06 $X=5735 $Y=20205 $D=2
M523 425 RDE vdd vdd p12ll L=6e-08 W=1.4e-06 $X=5745 $Y=9390 $D=2
M524 vdd vdd A[6] vdd p12ll L=6e-08 W=2e-07 $X=5810 $Y=5245 $D=2
M525 vdd 144 141 vdd p12ll L=6e-08 W=1.5e-06 $X=5860 $Y=15140 $D=2
M526 vdd 142 PXA[2] vdd p12ll L=6e-08 W=3.5e-06 $X=5880 $Y=26845 $D=2
M527 144 143 425 vdd p12ll L=6e-08 W=1.4e-06 $X=6035 $Y=9390 $D=2
M528 A[7] vdd vdd vdd p12ll L=6e-08 W=2e-07 $X=6090 $Y=5245 $D=2
M529 PXA[0] 146 vdd vdd p12ll L=6e-08 W=3.5e-06 $X=6220 $Y=26845 $D=2
M530 147 144 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=6240 $Y=15140 $D=2
M531 148 145 vdd vdd p12ll L=6e-08 W=4e-07 $X=6285 $Y=1395 $D=2
M532 149 PXA[1] vdd vdd p12ll L=3e-07 W=1.2e-07 $X=6315 $Y=31630 $D=2
M533 146 120 147 vdd p12ll L=6e-08 W=2.5e-06 $X=6365 $Y=20205 $D=2
M534 vdd 146 PXA[0] vdd p12ll L=6e-08 W=3.5e-06 $X=6510 $Y=26845 $D=2
M535 vdd 154 147 vdd p12ll L=6e-08 W=1.5e-06 $X=6520 $Y=15140 $D=2
M536 vdd PXA[0] 146 vdd p12ll L=3e-07 W=1.2e-07 $X=6570 $Y=30975 $D=2
M537 426 vss vdd vdd p12ll L=1e-07 W=4e-07 $X=6625 $Y=8465 $D=2
M538 151 154 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=6790 $Y=15140 $D=2
M539 PXA[1] 149 vdd vdd p12ll L=6e-08 W=3.5e-06 $X=6800 $Y=26845 $D=2
M540 vdd 153 150 vdd p12ll L=6e-08 W=1.4e-06 $X=6815 $Y=9390 $D=2
M541 vdd 148 155 vdd p12ll L=6e-08 W=1e-06 $X=6925 $Y=830 $D=2
M542 151 120 149 vdd p12ll L=6e-08 W=2.5e-06 $X=6945 $Y=20205 $D=2
M543 153 A[7] 426 vdd p12ll L=6e-08 W=4e-07 $X=6970 $Y=8465 $D=2
M544 vdd 152 151 vdd p12ll L=6e-08 W=1.5e-06 $X=7070 $Y=15140 $D=2
M545 vdd 149 PXA[1] vdd p12ll L=6e-08 W=3.5e-06 $X=7090 $Y=26845 $D=2
M546 154 150 vdd vdd p12ll L=6e-08 W=1.4e-06 $X=7105 $Y=9390 $D=2
M547 155 148 vdd vdd p12ll L=6e-08 W=1e-06 $X=7215 $Y=830 $D=2
M548 155 120 163 vdd p12ll L=6e-08 W=1.25e-06 $X=7875 $Y=580 $D=2
M549 163 120 155 vdd p12ll L=6e-08 W=1.25e-06 $X=8165 $Y=580 $D=2
M550 vdd vdd A[5] vdd p12ll L=6e-08 W=2e-07 $X=8580 $Y=13685 $D=2
M551 160 158 vdd vdd p12ll L=6e-08 W=4e-07 $X=8685 $Y=24100 $D=2
M552 FCKX[3] 158 180 vdd p12ll L=6e-08 W=1.25e-06 $X=8685 $Y=27295 $D=2
M553 FCKX[3] 160 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=8685 $Y=30855 $D=2
M554 161 120 158 vdd p12ll L=6e-08 W=5e-07 $X=8845 $Y=22145 $D=2
M555 A[3] vdd vdd vdd p12ll L=6e-08 W=2e-07 $X=8940 $Y=13685 $D=2
M556 vdd 159 161 vdd p12ll L=6e-08 W=1e-06 $X=8975 $Y=18030 $D=2
M557 vdd 158 160 vdd p12ll L=6e-08 W=4e-07 $X=8975 $Y=24100 $D=2
M558 180 158 FCKX[3] vdd p12ll L=6e-08 W=1.25e-06 $X=8975 $Y=27295 $D=2
M559 vdd 160 FCKX[3] vdd p12ll L=6e-08 W=1.25e-06 $X=8975 $Y=30855 $D=2
M560 158 120 161 vdd p12ll L=6e-08 W=5e-07 $X=9115 $Y=22145 $D=2
M561 vdd 160 158 vdd p12ll L=3e-07 W=1.2e-07 $X=9225 $Y=23260 $D=2
M562 161 162 vdd vdd p12ll L=6e-08 W=1e-06 $X=9265 $Y=18030 $D=2
M563 160 158 vdd vdd p12ll L=6e-08 W=4e-07 $X=9265 $Y=24100 $D=2
M564 FCKX[3] 158 180 vdd p12ll L=6e-08 W=1.25e-06 $X=9265 $Y=27295 $D=2
M565 FCKX[3] 160 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=9265 $Y=30855 $D=2
M566 161 120 158 vdd p12ll L=6e-08 W=5e-07 $X=9395 $Y=22145 $D=2
M567 174 199 vdd vdd p12ll L=6e-08 W=1e-06 $X=9465 $Y=16170 $D=2
M568 vdd 174 161 vdd p12ll L=6e-08 W=1e-06 $X=9555 $Y=18030 $D=2
M569 vdd 158 160 vdd p12ll L=6e-08 W=4e-07 $X=9555 $Y=24100 $D=2
M570 180 158 FCKX[3] vdd p12ll L=6e-08 W=1.25e-06 $X=9555 $Y=27295 $D=2
M571 vdd 160 FCKX[3] vdd p12ll L=6e-08 W=1.25e-06 $X=9555 $Y=30855 $D=2
M572 vdd 199 174 vdd p12ll L=6e-08 W=1e-06 $X=9755 $Y=16170 $D=2
M573 ZASX 163 vdd vdd p12ll L=6e-08 W=5.005e-06 $X=9815 $Y=8790 $D=2
M574 165 174 vdd vdd p12ll L=6e-08 W=1e-06 $X=9845 $Y=18030 $D=2
M575 164 166 vdd vdd p12ll L=6e-08 W=4e-07 $X=9845 $Y=24100 $D=2
M576 FCKX[2] 166 180 vdd p12ll L=6e-08 W=1.25e-06 $X=9845 $Y=27295 $D=2
M577 FCKX[2] 164 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=9845 $Y=30855 $D=2
M578 166 164 vdd vdd p12ll L=3e-07 W=1.2e-07 $X=9935 $Y=23260 $D=2
M579 166 120 165 vdd p12ll L=6e-08 W=5e-07 $X=10005 $Y=22145 $D=2
M580 199 168 vdd vdd p12ll L=6e-08 W=1e-06 $X=10045 $Y=16170 $D=2
M581 vdd ZASX 163 vdd p12ll L=3e-07 W=1.2e-07 $X=10095 $Y=1705 $D=2
M582 vdd 163 ZASX vdd p12ll L=6e-08 W=5.005e-06 $X=10105 $Y=8790 $D=2
M583 vdd 162 165 vdd p12ll L=6e-08 W=1e-06 $X=10135 $Y=18030 $D=2
M584 vdd 166 164 vdd p12ll L=6e-08 W=4e-07 $X=10135 $Y=24100 $D=2
M585 180 166 FCKX[2] vdd p12ll L=6e-08 W=1.25e-06 $X=10135 $Y=27295 $D=2
M586 vdd 164 FCKX[2] vdd p12ll L=6e-08 W=1.25e-06 $X=10135 $Y=30855 $D=2
M587 165 120 166 vdd p12ll L=6e-08 W=5e-07 $X=10285 $Y=22145 $D=2
M588 vdd 168 199 vdd p12ll L=6e-08 W=1e-06 $X=10335 $Y=16170 $D=2
M589 ZAS 170 vdd vdd p12ll L=6e-08 W=5.005e-06 $X=10395 $Y=8790 $D=2
M590 165 167 vdd vdd p12ll L=6e-08 W=1e-06 $X=10425 $Y=18030 $D=2
M591 164 166 vdd vdd p12ll L=6e-08 W=4e-07 $X=10425 $Y=24100 $D=2
M592 FCKX[2] 166 180 vdd p12ll L=6e-08 W=1.25e-06 $X=10425 $Y=27295 $D=2
M593 FCKX[2] 164 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=10425 $Y=30855 $D=2
M594 166 120 165 vdd p12ll L=6e-08 W=5e-07 $X=10555 $Y=22145 $D=2
M595 vdd 170 ZAS vdd p12ll L=6e-08 W=5.005e-06 $X=10685 $Y=8790 $D=2
M596 vdd 166 164 vdd p12ll L=6e-08 W=4e-07 $X=10715 $Y=24100 $D=2
M597 180 166 FCKX[2] vdd p12ll L=6e-08 W=1.25e-06 $X=10715 $Y=27295 $D=2
M598 vdd 164 FCKX[2] vdd p12ll L=6e-08 W=1.25e-06 $X=10715 $Y=30855 $D=2
M599 427 A[5] 168 vdd p12ll L=6e-08 W=4e-07 $X=10965 $Y=16500 $D=2
M600 172 169 vdd vdd p12ll L=6e-08 W=4e-07 $X=11005 $Y=24100 $D=2
M601 FCKX[0] 169 180 vdd p12ll L=6e-08 W=1.25e-06 $X=11005 $Y=27295 $D=2
M602 FCKX[0] 172 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=11005 $Y=30855 $D=2
M603 170 163 vdd vdd p12ll L=6e-08 W=2e-06 $X=11035 $Y=8790 $D=2
M604 171 CLK vdd vdd p12ll L=6e-08 W=4e-07 $X=11055 $Y=1620 $D=2
M605 CLK vdd vdd vdd p12ll L=6e-08 W=2e-07 $X=11140 $Y=765 $D=2
M606 173 120 169 vdd p12ll L=6e-08 W=5e-07 $X=11165 $Y=22145 $D=2
M607 vdd vss 427 vdd p12ll L=1e-07 W=4e-07 $X=11245 $Y=16500 $D=2
M608 vdd 167 173 vdd p12ll L=6e-08 W=1e-06 $X=11295 $Y=18030 $D=2
M609 vdd 169 172 vdd p12ll L=6e-08 W=4e-07 $X=11295 $Y=24100 $D=2
M610 180 169 FCKX[0] vdd p12ll L=6e-08 W=1.25e-06 $X=11295 $Y=27295 $D=2
M611 vdd 172 FCKX[0] vdd p12ll L=6e-08 W=1.25e-06 $X=11295 $Y=30855 $D=2
M612 169 120 173 vdd p12ll L=6e-08 W=5e-07 $X=11435 $Y=22145 $D=2
M613 vdd 172 169 vdd p12ll L=3e-07 W=1.2e-07 $X=11545 $Y=23260 $D=2
M614 173 207 vdd vdd p12ll L=6e-08 W=1e-06 $X=11585 $Y=18030 $D=2
M615 172 169 vdd vdd p12ll L=6e-08 W=4e-07 $X=11585 $Y=24100 $D=2
M616 FCKX[0] 169 180 vdd p12ll L=6e-08 W=1.25e-06 $X=11585 $Y=27295 $D=2
M617 FCKX[0] 172 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=11585 $Y=30855 $D=2
M618 173 120 169 vdd p12ll L=6e-08 W=5e-07 $X=11715 $Y=22145 $D=2
M619 vdd vdd CEN vdd p12ll L=6e-08 W=2e-07 $X=11735 $Y=1840 $D=2
M620 vdd 174 173 vdd p12ll L=6e-08 W=1e-06 $X=11875 $Y=18030 $D=2
M621 vdd 169 172 vdd p12ll L=6e-08 W=4e-07 $X=11875 $Y=24100 $D=2
M622 180 169 FCKX[0] vdd p12ll L=6e-08 W=1.25e-06 $X=11875 $Y=27295 $D=2
M623 vdd 172 FCKX[0] vdd p12ll L=6e-08 W=1.25e-06 $X=11875 $Y=30855 $D=2
M624 428 CLK vdd vdd p12ll L=6e-08 W=1e-06 $X=12075 $Y=1040 $D=2
M625 178 174 vdd vdd p12ll L=6e-08 W=1e-06 $X=12165 $Y=18030 $D=2
M626 176 177 vdd vdd p12ll L=6e-08 W=4e-07 $X=12165 $Y=24100 $D=2
M627 FCKX[1] 177 180 vdd p12ll L=6e-08 W=1.25e-06 $X=12165 $Y=27295 $D=2
M628 FCKX[1] 176 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=12165 $Y=30855 $D=2
M629 177 176 vdd vdd p12ll L=3e-07 W=1.2e-07 $X=12255 $Y=23260 $D=2
M630 175 CEN 428 vdd p12ll L=6e-08 W=1e-06 $X=12295 $Y=1040 $D=2
M631 177 120 178 vdd p12ll L=6e-08 W=5e-07 $X=12325 $Y=22145 $D=2
M632 181 179 vdd vdd p12ll L=6e-08 W=1.24e-06 $X=12330 $Y=11240 $D=2
M633 vdd 207 178 vdd p12ll L=6e-08 W=1e-06 $X=12455 $Y=18030 $D=2
M634 vdd 177 176 vdd p12ll L=6e-08 W=4e-07 $X=12455 $Y=24100 $D=2
M635 180 177 FCKX[1] vdd p12ll L=6e-08 W=1.25e-06 $X=12455 $Y=27295 $D=2
M636 vdd 176 FCKX[1] vdd p12ll L=6e-08 W=1.25e-06 $X=12455 $Y=30855 $D=2
M637 178 120 177 vdd p12ll L=6e-08 W=5e-07 $X=12605 $Y=22145 $D=2
M638 vdd 179 181 vdd p12ll L=6e-08 W=1.24e-06 $X=12620 $Y=11240 $D=2
M639 vdd 184 175 vdd p12ll L=3e-07 W=1.2e-07 $X=12650 $Y=1815 $D=2
M640 178 159 vdd vdd p12ll L=6e-08 W=1e-06 $X=12745 $Y=18030 $D=2
M641 176 177 vdd vdd p12ll L=6e-08 W=4e-07 $X=12745 $Y=24100 $D=2
M642 FCKX[1] 177 180 vdd p12ll L=6e-08 W=1.25e-06 $X=12745 $Y=27295 $D=2
M643 FCKX[1] 176 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=12745 $Y=30855 $D=2
M644 180 126 216 vdd p12ll L=6e-08 W=1e-06 $X=12810 $Y=33415 $D=2
M645 217 126 180 vdd p12ll L=6e-08 W=1e-06 $X=12810 $Y=33685 $D=2
M646 429 vss vdd vdd p12ll L=1e-07 W=4e-07 $X=12815 $Y=16500 $D=2
M647 177 120 178 vdd p12ll L=6e-08 W=5e-07 $X=12875 $Y=22145 $D=2
M648 179 DBL vdd vdd p12ll L=6e-08 W=8e-07 $X=12910 $Y=11680 $D=2
M649 vdd 177 176 vdd p12ll L=6e-08 W=4e-07 $X=13035 $Y=24100 $D=2
M650 180 177 FCKX[1] vdd p12ll L=6e-08 W=1.25e-06 $X=13035 $Y=27295 $D=2
M651 vdd 176 FCKX[1] vdd p12ll L=6e-08 W=1.25e-06 $X=13035 $Y=30855 $D=2
M652 183 A[3] 429 vdd p12ll L=6e-08 W=4e-07 $X=13135 $Y=16500 $D=2
M653 185 182 vdd vdd p12ll L=6e-08 W=4e-07 $X=13325 $Y=24100 $D=2
M654 FCKX[7] 182 180 vdd p12ll L=6e-08 W=1.25e-06 $X=13325 $Y=27295 $D=2
M655 FCKX[7] 185 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=13325 $Y=30855 $D=2
M656 186 120 182 vdd p12ll L=6e-08 W=5e-07 $X=13485 $Y=22145 $D=2
M657 vdd 175 184 vdd p12ll L=6e-08 W=8e-07 $X=13560 $Y=1240 $D=2
M658 vdd 159 186 vdd p12ll L=6e-08 W=1e-06 $X=13615 $Y=18030 $D=2
M659 vdd 182 185 vdd p12ll L=6e-08 W=4e-07 $X=13615 $Y=24100 $D=2
M660 180 182 FCKX[7] vdd p12ll L=6e-08 W=1.25e-06 $X=13615 $Y=27295 $D=2
M661 vdd 185 FCKX[7] vdd p12ll L=6e-08 W=1.25e-06 $X=13615 $Y=30855 $D=2
M662 EMCLK 187 vdd vdd p12ll L=6e-08 W=1.2e-06 $X=13690 $Y=11280 $D=2
M663 182 120 186 vdd p12ll L=6e-08 W=5e-07 $X=13755 $Y=22145 $D=2
M664 159 183 vdd vdd p12ll L=6e-08 W=1e-06 $X=13765 $Y=16170 $D=2
M665 DBL 201 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=13835 $Y=9085 $D=2
M666 430 184 vdd vdd p12ll L=6e-08 W=1e-06 $X=13850 $Y=1040 $D=2
M667 vdd 185 182 vdd p12ll L=3e-07 W=1.2e-07 $X=13865 $Y=23260 $D=2
M668 186 162 vdd vdd p12ll L=6e-08 W=1e-06 $X=13905 $Y=18030 $D=2
M669 185 182 vdd vdd p12ll L=6e-08 W=4e-07 $X=13905 $Y=24100 $D=2
M670 FCKX[7] 182 180 vdd p12ll L=6e-08 W=1.25e-06 $X=13905 $Y=27295 $D=2
M671 FCKX[7] 185 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=13905 $Y=30855 $D=2
M672 vdd 187 EMCLK vdd p12ll L=6e-08 W=1.2e-06 $X=13980 $Y=11280 $D=2
M673 186 120 182 vdd p12ll L=6e-08 W=5e-07 $X=14035 $Y=22145 $D=2
M674 vdd 183 159 vdd p12ll L=6e-08 W=1e-06 $X=14055 $Y=16170 $D=2
M675 vdd 201 DBL vdd p12ll L=6e-08 W=1.25e-06 $X=14125 $Y=9085 $D=2
M676 188 CLK 430 vdd p12ll L=6e-08 W=1e-06 $X=14140 $Y=1040 $D=2
M677 vdd 199 186 vdd p12ll L=6e-08 W=1e-06 $X=14195 $Y=18030 $D=2
M678 vdd 182 185 vdd p12ll L=6e-08 W=4e-07 $X=14195 $Y=24100 $D=2
M679 180 182 FCKX[7] vdd p12ll L=6e-08 W=1.25e-06 $X=14195 $Y=27295 $D=2
M680 vdd 185 FCKX[7] vdd p12ll L=6e-08 W=1.25e-06 $X=14195 $Y=30855 $D=2
M681 167 159 vdd vdd p12ll L=6e-08 W=1e-06 $X=14345 $Y=16170 $D=2
M682 202 181 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=14415 $Y=9085 $D=2
M683 190 199 vdd vdd p12ll L=6e-08 W=1e-06 $X=14485 $Y=18030 $D=2
M684 189 191 vdd vdd p12ll L=6e-08 W=4e-07 $X=14485 $Y=24100 $D=2
M685 FCKX[6] 191 180 vdd p12ll L=6e-08 W=1.25e-06 $X=14485 $Y=27295 $D=2
M686 FCKX[6] 189 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=14485 $Y=30855 $D=2
M687 191 189 vdd vdd p12ll L=3e-07 W=1.2e-07 $X=14575 $Y=23260 $D=2
M688 vdd 159 167 vdd p12ll L=6e-08 W=1e-06 $X=14635 $Y=16170 $D=2
M689 191 120 190 vdd p12ll L=6e-08 W=5e-07 $X=14645 $Y=22145 $D=2
M690 vdd 181 202 vdd p12ll L=6e-08 W=1.25e-06 $X=14705 $Y=9085 $D=2
M691 vdd 192 187 vdd p12ll L=6e-08 W=6e-07 $X=14745 $Y=11880 $D=2
M692 vdd 162 190 vdd p12ll L=6e-08 W=1e-06 $X=14775 $Y=18030 $D=2
M693 vdd 191 189 vdd p12ll L=6e-08 W=4e-07 $X=14775 $Y=24100 $D=2
M694 180 191 FCKX[6] vdd p12ll L=6e-08 W=1.25e-06 $X=14775 $Y=27295 $D=2
M695 vdd 189 FCKX[6] vdd p12ll L=6e-08 W=1.25e-06 $X=14775 $Y=30855 $D=2
M696 vdd 188 193 vdd p12ll L=6e-08 W=1e-06 $X=14830 $Y=1170 $D=2
M697 190 120 191 vdd p12ll L=6e-08 W=5e-07 $X=14925 $Y=22145 $D=2
M698 202 181 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=14995 $Y=9085 $D=2
M699 192 197 vdd vdd p12ll L=6e-08 W=6e-07 $X=15035 $Y=11880 $D=2
M700 190 167 vdd vdd p12ll L=6e-08 W=1e-06 $X=15065 $Y=18030 $D=2
M701 189 191 vdd vdd p12ll L=6e-08 W=4e-07 $X=15065 $Y=24100 $D=2
M702 FCKX[6] 191 180 vdd p12ll L=6e-08 W=1.25e-06 $X=15065 $Y=27295 $D=2
M703 FCKX[6] 189 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=15065 $Y=30855 $D=2
M704 194 193 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=15180 $Y=670 $D=2
M705 191 120 190 vdd p12ll L=6e-08 W=5e-07 $X=15195 $Y=22145 $D=2
M706 vdd 181 202 vdd p12ll L=6e-08 W=1.25e-06 $X=15285 $Y=9085 $D=2
M707 vdd 191 189 vdd p12ll L=6e-08 W=4e-07 $X=15355 $Y=24100 $D=2
M708 180 191 FCKX[6] vdd p12ll L=6e-08 W=1.25e-06 $X=15355 $Y=27295 $D=2
M709 vdd 189 FCKX[6] vdd p12ll L=6e-08 W=1.25e-06 $X=15355 $Y=30855 $D=2
M710 vdd 193 194 vdd p12ll L=6e-08 W=1.5e-06 $X=15470 $Y=670 $D=2
M711 202 181 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=15575 $Y=9085 $D=2
M712 196 195 vdd vdd p12ll L=6e-08 W=4e-07 $X=15645 $Y=24100 $D=2
M713 FCKX[4] 195 180 vdd p12ll L=6e-08 W=1.25e-06 $X=15645 $Y=27295 $D=2
M714 FCKX[4] 196 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=15645 $Y=30855 $D=2
M715 431 vss vdd vdd p12ll L=1e-07 W=4e-07 $X=15715 $Y=16500 $D=2
M716 198 120 195 vdd p12ll L=6e-08 W=5e-07 $X=15805 $Y=22145 $D=2
M717 vdd 181 202 vdd p12ll L=6e-08 W=1.25e-06 $X=15865 $Y=9085 $D=2
M718 221 215 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=15870 $Y=670 $D=2
M719 vdd 167 198 vdd p12ll L=6e-08 W=1e-06 $X=15935 $Y=18030 $D=2
M720 vdd 195 196 vdd p12ll L=6e-08 W=4e-07 $X=15935 $Y=24100 $D=2
M721 180 195 FCKX[4] vdd p12ll L=6e-08 W=1.25e-06 $X=15935 $Y=27295 $D=2
M722 vdd 196 FCKX[4] vdd p12ll L=6e-08 W=1.25e-06 $X=15935 $Y=30855 $D=2
M723 200 A[4] 431 vdd p12ll L=6e-08 W=4e-07 $X=16035 $Y=16500 $D=2
M724 vdd 129 216 vdd p12ll L=6e-08 W=2e-06 $X=16065 $Y=33415 $D=2
M725 217 129 vdd vdd p12ll L=6e-08 W=2e-06 $X=16065 $Y=33685 $D=2
M726 195 120 198 vdd p12ll L=6e-08 W=5e-07 $X=16075 $Y=22145 $D=2
M727 202 181 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=16155 $Y=9085 $D=2
M728 vdd 215 221 vdd p12ll L=6e-08 W=1.5e-06 $X=16185 $Y=670 $D=2
M729 vdd 196 195 vdd p12ll L=3e-07 W=1.2e-07 $X=16185 $Y=23260 $D=2
M730 198 207 vdd vdd p12ll L=6e-08 W=1e-06 $X=16225 $Y=18030 $D=2
M731 196 195 vdd vdd p12ll L=6e-08 W=4e-07 $X=16225 $Y=24100 $D=2
M732 FCKX[4] 195 180 vdd p12ll L=6e-08 W=1.25e-06 $X=16225 $Y=27295 $D=2
M733 FCKX[4] 196 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=16225 $Y=30855 $D=2
M734 vdd 201 197 vdd p12ll L=6e-08 W=6e-07 $X=16320 $Y=11880 $D=2
M735 198 120 195 vdd p12ll L=6e-08 W=5e-07 $X=16355 $Y=22145 $D=2
M736 vdd 181 202 vdd p12ll L=6e-08 W=1.25e-06 $X=16445 $Y=9085 $D=2
M737 vdd 199 198 vdd p12ll L=6e-08 W=1e-06 $X=16515 $Y=18030 $D=2
M738 vdd 195 196 vdd p12ll L=6e-08 W=4e-07 $X=16515 $Y=24100 $D=2
M739 180 195 FCKX[4] vdd p12ll L=6e-08 W=1.25e-06 $X=16515 $Y=27295 $D=2
M740 vdd 196 FCKX[4] vdd p12ll L=6e-08 W=1.25e-06 $X=16515 $Y=30855 $D=2
M741 203 251 vdd vdd p12ll L=6e-08 W=1.5e-06 $X=16540 $Y=670 $D=2
M742 162 200 vdd vdd p12ll L=6e-08 W=1e-06 $X=16665 $Y=16170 $D=2
M743 201 202 vdd vdd p12ll L=6e-08 W=1.4e-06 $X=16670 $Y=11080 $D=2
M744 210 199 vdd vdd p12ll L=6e-08 W=1e-06 $X=16805 $Y=18030 $D=2
M745 206 208 vdd vdd p12ll L=6e-08 W=4e-07 $X=16805 $Y=24100 $D=2
M746 FCKX[5] 208 180 vdd p12ll L=6e-08 W=1.25e-06 $X=16805 $Y=27295 $D=2
M747 FCKX[5] 206 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=16805 $Y=30855 $D=2
M748 204 211 203 vdd p12ll L=6e-08 W=1.5e-06 $X=16830 $Y=670 $D=2
M749 208 206 vdd vdd p12ll L=3e-07 W=1.2e-07 $X=16895 $Y=23260 $D=2
M750 vdd 200 162 vdd p12ll L=6e-08 W=1e-06 $X=16955 $Y=16170 $D=2
M751 208 120 210 vdd p12ll L=6e-08 W=5e-07 $X=16965 $Y=22145 $D=2
M752 vdd 207 210 vdd p12ll L=6e-08 W=1e-06 $X=17095 $Y=18030 $D=2
M753 vdd 208 206 vdd p12ll L=6e-08 W=4e-07 $X=17095 $Y=24100 $D=2
M754 180 208 FCKX[5] vdd p12ll L=6e-08 W=1.25e-06 $X=17095 $Y=27295 $D=2
M755 vdd 206 FCKX[5] vdd p12ll L=6e-08 W=1.25e-06 $X=17095 $Y=30855 $D=2
M756 203 211 204 vdd p12ll L=6e-08 W=1.5e-06 $X=17120 $Y=670 $D=2
M757 207 162 vdd vdd p12ll L=6e-08 W=1e-06 $X=17245 $Y=16170 $D=2
M758 210 120 208 vdd p12ll L=6e-08 W=5e-07 $X=17245 $Y=22145 $D=2
M759 210 159 vdd vdd p12ll L=6e-08 W=1e-06 $X=17385 $Y=18030 $D=2
M760 206 208 vdd vdd p12ll L=6e-08 W=4e-07 $X=17385 $Y=24100 $D=2
M761 FCKX[5] 208 180 vdd p12ll L=6e-08 W=1.25e-06 $X=17385 $Y=27295 $D=2
M762 FCKX[5] 206 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=17385 $Y=30855 $D=2
M763 vdd 251 203 vdd p12ll L=6e-08 W=1.5e-06 $X=17410 $Y=670 $D=2
M764 208 120 210 vdd p12ll L=6e-08 W=5e-07 $X=17515 $Y=22145 $D=2
M765 vdd 162 207 vdd p12ll L=6e-08 W=1e-06 $X=17535 $Y=16170 $D=2
M766 vdd 208 206 vdd p12ll L=6e-08 W=4e-07 $X=17675 $Y=24100 $D=2
M767 180 208 FCKX[5] vdd p12ll L=6e-08 W=1.25e-06 $X=17675 $Y=27295 $D=2
M768 vdd 206 FCKX[5] vdd p12ll L=6e-08 W=1.25e-06 $X=17675 $Y=30855 $D=2
M769 432 209 215 vdd p12ll L=6e-08 W=2.5e-06 $X=17760 $Y=8735 $D=2
M770 vdd vdd A[4] vdd p12ll L=6e-08 W=2e-07 $X=17955 $Y=14135 $D=2
M771 214 212 vdd vdd p12ll L=6e-08 W=4e-07 $X=17965 $Y=24100 $D=2
M772 YX[3] 212 180 vdd p12ll L=6e-08 W=1.25e-06 $X=17965 $Y=27295 $D=2
M773 YX[3] 214 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=17965 $Y=30855 $D=2
M774 vdd 251 432 vdd p12ll L=6e-08 W=2.5e-06 $X=18000 $Y=8735 $D=2
M775 vdd 219 211 vdd p12ll L=2e-07 W=4e-07 $X=18100 $Y=1465 $D=2
M776 218 120 212 vdd p12ll L=6e-08 W=5e-07 $X=18125 $Y=22145 $D=2
M777 vdd 213 218 vdd p12ll L=6e-08 W=1e-06 $X=18255 $Y=18030 $D=2
M778 vdd 212 214 vdd p12ll L=6e-08 W=4e-07 $X=18255 $Y=24100 $D=2
M779 180 212 YX[3] vdd p12ll L=6e-08 W=1.25e-06 $X=18255 $Y=27295 $D=2
M780 vdd 214 YX[3] vdd p12ll L=6e-08 W=1.25e-06 $X=18255 $Y=30855 $D=2
M781 A[2] vdd vdd vdd p12ll L=6e-08 W=2e-07 $X=18305 $Y=14135 $D=2
M782 120 215 vdd vdd p12ll L=6e-08 W=5e-06 $X=18340 $Y=8735 $D=2
M783 212 120 218 vdd p12ll L=6e-08 W=5e-07 $X=18395 $Y=22145 $D=2
M784 vdd 214 212 vdd p12ll L=3e-07 W=1.2e-07 $X=18505 $Y=23260 $D=2
M785 218 220 vdd vdd p12ll L=6e-08 W=1e-06 $X=18545 $Y=18030 $D=2
M786 214 212 vdd vdd p12ll L=6e-08 W=4e-07 $X=18545 $Y=24100 $D=2
M787 YX[3] 212 180 vdd p12ll L=6e-08 W=1.25e-06 $X=18545 $Y=27295 $D=2
M788 YX[3] 214 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=18545 $Y=30855 $D=2
M789 202 251 vdd vdd p12ll L=2e-07 W=1.2e-07 $X=18590 $Y=947 $D=2
M790 219 251 vdd vdd p12ll L=2e-07 W=4e-07 $X=18590 $Y=1465 $D=2
M791 vdd 215 120 vdd p12ll L=6e-08 W=5e-06 $X=18630 $Y=8735 $D=2
M792 218 120 212 vdd p12ll L=6e-08 W=5e-07 $X=18675 $Y=22145 $D=2
M793 231 249 vdd vdd p12ll L=6e-08 W=1e-06 $X=18745 $Y=16170 $D=2
M794 vdd 231 218 vdd p12ll L=6e-08 W=1e-06 $X=18835 $Y=18030 $D=2
M795 vdd 212 214 vdd p12ll L=6e-08 W=4e-07 $X=18835 $Y=24100 $D=2
M796 180 212 YX[3] vdd p12ll L=6e-08 W=1.25e-06 $X=18835 $Y=27295 $D=2
M797 vdd 214 YX[3] vdd p12ll L=6e-08 W=1.25e-06 $X=18835 $Y=30855 $D=2
M798 DCTRCLK 215 vdd vdd p12ll L=6e-08 W=5e-06 $X=18920 $Y=8735 $D=2
M799 vdd 249 231 vdd p12ll L=6e-08 W=1e-06 $X=19035 $Y=16170 $D=2
M800 223 231 vdd vdd p12ll L=6e-08 W=1e-06 $X=19125 $Y=18030 $D=2
M801 222 224 vdd vdd p12ll L=6e-08 W=4e-07 $X=19125 $Y=24100 $D=2
M802 YX[2] 224 180 vdd p12ll L=6e-08 W=1.25e-06 $X=19125 $Y=27295 $D=2
M803 YX[2] 222 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=19125 $Y=30855 $D=2
M804 vdd 215 DCTRCLK vdd p12ll L=6e-08 W=5e-06 $X=19210 $Y=8735 $D=2
M805 224 222 vdd vdd p12ll L=3e-07 W=1.2e-07 $X=19215 $Y=23260 $D=2
M806 224 120 223 vdd p12ll L=6e-08 W=5e-07 $X=19285 $Y=22145 $D=2
M807 249 226 vdd vdd p12ll L=6e-08 W=1e-06 $X=19325 $Y=16170 $D=2
M808 vdd 228 209 vdd p12ll L=2e-07 W=4e-07 $X=19410 $Y=1465 $D=2
M809 vdd 220 223 vdd p12ll L=6e-08 W=1e-06 $X=19415 $Y=18030 $D=2
M810 vdd 224 222 vdd p12ll L=6e-08 W=4e-07 $X=19415 $Y=24100 $D=2
M811 180 224 YX[2] vdd p12ll L=6e-08 W=1.25e-06 $X=19415 $Y=27295 $D=2
M812 vdd 222 YX[2] vdd p12ll L=6e-08 W=1.25e-06 $X=19415 $Y=30855 $D=2
M813 121 120 vdd vdd p12ll L=6e-08 W=5e-06 $X=19500 $Y=8735 $D=2
M814 223 120 224 vdd p12ll L=6e-08 W=5e-07 $X=19565 $Y=22145 $D=2
M815 vdd 226 249 vdd p12ll L=6e-08 W=1e-06 $X=19615 $Y=16170 $D=2
M816 223 225 vdd vdd p12ll L=6e-08 W=1e-06 $X=19705 $Y=18030 $D=2
M817 222 224 vdd vdd p12ll L=6e-08 W=4e-07 $X=19705 $Y=24100 $D=2
M818 YX[2] 224 180 vdd p12ll L=6e-08 W=1.25e-06 $X=19705 $Y=27295 $D=2
M819 YX[2] 222 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=19705 $Y=30855 $D=2
M820 vdd 120 121 vdd p12ll L=6e-08 W=5e-06 $X=19790 $Y=8735 $D=2
M821 224 120 223 vdd p12ll L=6e-08 W=5e-07 $X=19835 $Y=22145 $D=2
M822 433 vss vdd vdd p12ll L=2e-07 W=8e-07 $X=19900 $Y=1065 $D=2
M823 vdd 224 222 vdd p12ll L=6e-08 W=4e-07 $X=19995 $Y=24100 $D=2
M824 180 224 YX[2] vdd p12ll L=6e-08 W=1.25e-06 $X=19995 $Y=27295 $D=2
M825 vdd 222 YX[2] vdd p12ll L=6e-08 W=1.25e-06 $X=19995 $Y=30855 $D=2
M826 DCTRCLKX 221 vdd vdd p12ll L=6e-08 W=5e-06 $X=20080 $Y=8735 $D=2
M827 434 A[2] 226 vdd p12ll L=6e-08 W=4e-07 $X=20245 $Y=16500 $D=2
M828 229 227 vdd vdd p12ll L=6e-08 W=4e-07 $X=20285 $Y=24100 $D=2
M829 YX[0] 227 180 vdd p12ll L=6e-08 W=1.25e-06 $X=20285 $Y=27295 $D=2
M830 YX[0] 229 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=20285 $Y=30855 $D=2
M831 vdd 221 DCTRCLKX vdd p12ll L=6e-08 W=5e-06 $X=20370 $Y=8735 $D=2
M832 228 251 433 vdd p12ll L=2e-07 W=8e-07 $X=20390 $Y=1065 $D=2
M833 230 120 227 vdd p12ll L=6e-08 W=5e-07 $X=20445 $Y=22145 $D=2
M834 vdd vss 434 vdd p12ll L=1e-07 W=4e-07 $X=20525 $Y=16500 $D=2
M835 vdd 225 230 vdd p12ll L=6e-08 W=1e-06 $X=20575 $Y=18030 $D=2
M836 vdd 227 229 vdd p12ll L=6e-08 W=4e-07 $X=20575 $Y=24100 $D=2
M837 180 227 YX[0] vdd p12ll L=6e-08 W=1.25e-06 $X=20575 $Y=27295 $D=2
M838 vdd 229 YX[0] vdd p12ll L=6e-08 W=1.25e-06 $X=20575 $Y=30855 $D=2
M839 SACK4 204 vdd vdd p12ll L=6e-08 W=5e-06 $X=20660 $Y=8735 $D=2
M840 227 120 230 vdd p12ll L=6e-08 W=5e-07 $X=20715 $Y=22145 $D=2
M841 vdd 229 227 vdd p12ll L=3e-07 W=1.2e-07 $X=20825 $Y=23260 $D=2
M842 230 254 vdd vdd p12ll L=6e-08 W=1e-06 $X=20865 $Y=18030 $D=2
M843 229 227 vdd vdd p12ll L=6e-08 W=4e-07 $X=20865 $Y=24100 $D=2
M844 YX[0] 227 180 vdd p12ll L=6e-08 W=1.25e-06 $X=20865 $Y=27295 $D=2
M845 YX[0] 229 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=20865 $Y=30855 $D=2
M846 vdd 204 SACK4 vdd p12ll L=6e-08 W=5e-06 $X=20950 $Y=8735 $D=2
M847 230 120 227 vdd p12ll L=6e-08 W=5e-07 $X=20995 $Y=22145 $D=2
M848 WEN vdd vdd vdd p12ll L=6e-08 W=2e-07 $X=21055 $Y=490 $D=2
M849 vdd 231 230 vdd p12ll L=6e-08 W=1e-06 $X=21155 $Y=18030 $D=2
M850 vdd 227 229 vdd p12ll L=6e-08 W=4e-07 $X=21155 $Y=24100 $D=2
M851 180 227 YX[0] vdd p12ll L=6e-08 W=1.25e-06 $X=21155 $Y=27295 $D=2
M852 vdd 229 YX[0] vdd p12ll L=6e-08 W=1.25e-06 $X=21155 $Y=30855 $D=2
M853 vdd WEN 232 vdd p12ll L=6e-08 W=4e-07 $X=21180 $Y=1565 $D=2
M854 251 202 vdd vdd p12ll L=6e-08 W=5e-06 $X=21240 $Y=8735 $D=2
M855 vdd 216 RWLL vdd p12ll L=6e-08 W=5e-06 $X=21365 $Y=33415 $D=2
M856 RWLR 217 vdd vdd p12ll L=6e-08 W=5e-06 $X=21365 $Y=33685 $D=2
M857 235 231 vdd vdd p12ll L=6e-08 W=1e-06 $X=21445 $Y=18030 $D=2
M858 233 234 vdd vdd p12ll L=6e-08 W=4e-07 $X=21445 $Y=24100 $D=2
M859 YX[1] 234 180 vdd p12ll L=6e-08 W=1.25e-06 $X=21445 $Y=27295 $D=2
M860 YX[1] 233 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=21445 $Y=30855 $D=2
M861 236 232 vdd vdd p12ll L=3e-07 W=4e-07 $X=21500 $Y=1565 $D=2
M862 vdd 202 251 vdd p12ll L=6e-08 W=5e-06 $X=21530 $Y=8735 $D=2
M863 234 233 vdd vdd p12ll L=3e-07 W=1.2e-07 $X=21535 $Y=23260 $D=2
M864 234 120 235 vdd p12ll L=6e-08 W=5e-07 $X=21605 $Y=22145 $D=2
M865 vdd 254 235 vdd p12ll L=6e-08 W=1e-06 $X=21735 $Y=18030 $D=2
M866 vdd 234 233 vdd p12ll L=6e-08 W=4e-07 $X=21735 $Y=24100 $D=2
M867 180 234 YX[1] vdd p12ll L=6e-08 W=1.25e-06 $X=21735 $Y=27295 $D=2
M868 vdd 233 YX[1] vdd p12ll L=6e-08 W=1.25e-06 $X=21735 $Y=30855 $D=2
M869 251 202 vdd vdd p12ll L=6e-08 W=5e-06 $X=21820 $Y=8735 $D=2
M870 235 120 234 vdd p12ll L=6e-08 W=5e-07 $X=21885 $Y=22145 $D=2
M871 235 213 vdd vdd p12ll L=6e-08 W=1e-06 $X=22025 $Y=18030 $D=2
M872 233 234 vdd vdd p12ll L=6e-08 W=4e-07 $X=22025 $Y=24100 $D=2
M873 YX[1] 234 180 vdd p12ll L=6e-08 W=1.25e-06 $X=22025 $Y=27295 $D=2
M874 YX[1] 233 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=22025 $Y=30855 $D=2
M875 435 vss vdd vdd p12ll L=1e-07 W=4e-07 $X=22095 $Y=16500 $D=2
M876 vdd 202 251 vdd p12ll L=6e-08 W=5e-06 $X=22110 $Y=8735 $D=2
M877 234 120 235 vdd p12ll L=6e-08 W=5e-07 $X=22155 $Y=22145 $D=2
M878 vdd 234 233 vdd p12ll L=6e-08 W=4e-07 $X=22315 $Y=24100 $D=2
M879 180 234 YX[1] vdd p12ll L=6e-08 W=1.25e-06 $X=22315 $Y=27295 $D=2
M880 vdd 233 YX[1] vdd p12ll L=6e-08 W=1.25e-06 $X=22315 $Y=30855 $D=2
M881 SACK1 251 vdd vdd p12ll L=6e-08 W=5e-06 $X=22400 $Y=8735 $D=2
M882 238 A[0] 435 vdd p12ll L=6e-08 W=4e-07 $X=22415 $Y=16500 $D=2
M883 vdd 236 239 vdd p12ll L=2e-07 W=4e-07 $X=22460 $Y=1565 $D=2
M884 241 237 vdd vdd p12ll L=6e-08 W=4e-07 $X=22605 $Y=24100 $D=2
M885 YX[7] 237 180 vdd p12ll L=6e-08 W=1.25e-06 $X=22605 $Y=27295 $D=2
M886 YX[7] 241 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=22605 $Y=30855 $D=2
M887 vdd 251 SACK1 vdd p12ll L=6e-08 W=5e-06 $X=22690 $Y=8735 $D=2
M888 242 120 237 vdd p12ll L=6e-08 W=5e-07 $X=22765 $Y=22145 $D=2
M889 vdd 213 242 vdd p12ll L=6e-08 W=1e-06 $X=22895 $Y=18030 $D=2
M890 vdd 237 241 vdd p12ll L=6e-08 W=4e-07 $X=22895 $Y=24100 $D=2
M891 180 237 YX[7] vdd p12ll L=6e-08 W=1.25e-06 $X=22895 $Y=27295 $D=2
M892 vdd 241 YX[7] vdd p12ll L=6e-08 W=1.25e-06 $X=22895 $Y=30855 $D=2
M893 180 251 vdd vdd p12ll L=6e-08 W=2.5e-06 $X=22980 $Y=8735 $D=2
M894 240 239 vdd vdd p12ll L=6e-08 W=1e-06 $X=22995 $Y=965 $D=2
M895 237 120 242 vdd p12ll L=6e-08 W=5e-07 $X=23035 $Y=22145 $D=2
M896 213 238 vdd vdd p12ll L=6e-08 W=1e-06 $X=23045 $Y=16170 $D=2
M897 vdd 241 237 vdd p12ll L=3e-07 W=1.2e-07 $X=23145 $Y=23260 $D=2
M898 242 220 vdd vdd p12ll L=6e-08 W=1e-06 $X=23185 $Y=18030 $D=2
M899 241 237 vdd vdd p12ll L=6e-08 W=4e-07 $X=23185 $Y=24100 $D=2
M900 YX[7] 237 180 vdd p12ll L=6e-08 W=1.25e-06 $X=23185 $Y=27295 $D=2
M901 YX[7] 241 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=23185 $Y=30855 $D=2
M902 vdd 251 180 vdd p12ll L=6e-08 W=2.5e-06 $X=23270 $Y=8735 $D=2
M903 257 120 240 vdd p12ll L=6e-08 W=1e-06 $X=23285 $Y=965 $D=2
M904 242 120 237 vdd p12ll L=6e-08 W=5e-07 $X=23315 $Y=22145 $D=2
M905 vdd 238 213 vdd p12ll L=6e-08 W=1e-06 $X=23335 $Y=16170 $D=2
M906 vdd 249 242 vdd p12ll L=6e-08 W=1e-06 $X=23475 $Y=18030 $D=2
M907 vdd 237 241 vdd p12ll L=6e-08 W=4e-07 $X=23475 $Y=24100 $D=2
M908 180 237 YX[7] vdd p12ll L=6e-08 W=1.25e-06 $X=23475 $Y=27295 $D=2
M909 vdd 241 YX[7] vdd p12ll L=6e-08 W=1.25e-06 $X=23475 $Y=30855 $D=2
M910 180 251 vdd vdd p12ll L=6e-08 W=2.5e-06 $X=23560 $Y=8735 $D=2
M911 225 213 vdd vdd p12ll L=6e-08 W=1e-06 $X=23625 $Y=16170 $D=2
M912 244 249 vdd vdd p12ll L=6e-08 W=1e-06 $X=23765 $Y=18030 $D=2
M913 243 245 vdd vdd p12ll L=6e-08 W=4e-07 $X=23765 $Y=24100 $D=2
M914 YX[6] 245 180 vdd p12ll L=6e-08 W=1.25e-06 $X=23765 $Y=27295 $D=2
M915 YX[6] 243 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=23765 $Y=30855 $D=2
M916 vdd 251 180 vdd p12ll L=6e-08 W=2.5e-06 $X=23850 $Y=8735 $D=2
M917 245 243 vdd vdd p12ll L=3e-07 W=1.2e-07 $X=23855 $Y=23260 $D=2
M918 vdd 213 225 vdd p12ll L=6e-08 W=1e-06 $X=23915 $Y=16170 $D=2
M919 245 120 244 vdd p12ll L=6e-08 W=5e-07 $X=23925 $Y=22145 $D=2
M920 vdd vdd A[0] vdd p12ll L=6e-08 W=2e-07 $X=24025 $Y=1500 $D=2
M921 vdd 220 244 vdd p12ll L=6e-08 W=1e-06 $X=24055 $Y=18030 $D=2
M922 vdd 245 243 vdd p12ll L=6e-08 W=4e-07 $X=24055 $Y=24100 $D=2
M923 180 245 YX[6] vdd p12ll L=6e-08 W=1.25e-06 $X=24055 $Y=27295 $D=2
M924 vdd 243 YX[6] vdd p12ll L=6e-08 W=1.25e-06 $X=24055 $Y=30855 $D=2
M925 244 120 245 vdd p12ll L=6e-08 W=5e-07 $X=24205 $Y=22145 $D=2
M926 244 225 vdd vdd p12ll L=6e-08 W=1e-06 $X=24345 $Y=18030 $D=2
M927 243 245 vdd vdd p12ll L=6e-08 W=4e-07 $X=24345 $Y=24100 $D=2
M928 YX[6] 245 180 vdd p12ll L=6e-08 W=1.25e-06 $X=24345 $Y=27295 $D=2
M929 YX[6] 243 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=24345 $Y=30855 $D=2
M930 245 120 244 vdd p12ll L=6e-08 W=5e-07 $X=24475 $Y=22145 $D=2
M931 vdd 245 243 vdd p12ll L=6e-08 W=4e-07 $X=24635 $Y=24100 $D=2
M932 180 245 YX[6] vdd p12ll L=6e-08 W=1.25e-06 $X=24635 $Y=27295 $D=2
M933 vdd 243 YX[6] vdd p12ll L=6e-08 W=1.25e-06 $X=24635 $Y=30855 $D=2
M934 247 246 vdd vdd p12ll L=6e-08 W=4e-07 $X=24925 $Y=24100 $D=2
M935 YX[4] 246 180 vdd p12ll L=6e-08 W=1.25e-06 $X=24925 $Y=27295 $D=2
M936 YX[4] 247 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=24925 $Y=30855 $D=2
M937 436 vss vdd vdd p12ll L=1e-07 W=4e-07 $X=24995 $Y=16500 $D=2
M938 248 120 246 vdd p12ll L=6e-08 W=5e-07 $X=25085 $Y=22145 $D=2
M939 vdd 225 248 vdd p12ll L=6e-08 W=1e-06 $X=25215 $Y=18030 $D=2
M940 vdd 246 247 vdd p12ll L=6e-08 W=4e-07 $X=25215 $Y=24100 $D=2
M941 180 246 YX[4] vdd p12ll L=6e-08 W=1.25e-06 $X=25215 $Y=27295 $D=2
M942 vdd 247 YX[4] vdd p12ll L=6e-08 W=1.25e-06 $X=25215 $Y=30855 $D=2
M943 WE 252 vdd vdd p12ll L=6e-08 W=5e-06 $X=25300 $Y=8735 $D=2
M944 250 A[1] 436 vdd p12ll L=6e-08 W=4e-07 $X=25315 $Y=16500 $D=2
M945 246 120 248 vdd p12ll L=6e-08 W=5e-07 $X=25355 $Y=22145 $D=2
M946 vdd 247 246 vdd p12ll L=3e-07 W=1.2e-07 $X=25465 $Y=23260 $D=2
M947 248 254 vdd vdd p12ll L=6e-08 W=1e-06 $X=25505 $Y=18030 $D=2
M948 247 246 vdd vdd p12ll L=6e-08 W=4e-07 $X=25505 $Y=24100 $D=2
M949 YX[4] 246 180 vdd p12ll L=6e-08 W=1.25e-06 $X=25505 $Y=27295 $D=2
M950 YX[4] 247 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=25505 $Y=30855 $D=2
M951 vdd 252 WE vdd p12ll L=6e-08 W=5e-06 $X=25590 $Y=8735 $D=2
M952 248 120 246 vdd p12ll L=6e-08 W=5e-07 $X=25635 $Y=22145 $D=2
M953 vdd 249 248 vdd p12ll L=6e-08 W=1e-06 $X=25795 $Y=18030 $D=2
M954 vdd 246 247 vdd p12ll L=6e-08 W=4e-07 $X=25795 $Y=24100 $D=2
M955 180 246 YX[4] vdd p12ll L=6e-08 W=1.25e-06 $X=25795 $Y=27295 $D=2
M956 vdd 247 YX[4] vdd p12ll L=6e-08 W=1.25e-06 $X=25795 $Y=30855 $D=2
M957 vdd vdd A[1] vdd p12ll L=6e-08 W=2e-07 $X=25820 $Y=13980 $D=2
M958 252 258 vdd vdd p12ll L=6e-08 W=2.995e-06 $X=25880 $Y=8735 $D=2
M959 220 250 vdd vdd p12ll L=6e-08 W=1e-06 $X=25945 $Y=16170 $D=2
M960 256 249 vdd vdd p12ll L=6e-08 W=1e-06 $X=26085 $Y=18030 $D=2
M961 253 255 vdd vdd p12ll L=6e-08 W=4e-07 $X=26085 $Y=24100 $D=2
M962 YX[5] 255 180 vdd p12ll L=6e-08 W=1.25e-06 $X=26085 $Y=27295 $D=2
M963 YX[5] 253 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=26085 $Y=30855 $D=2
M964 vdd 251 252 vdd p12ll L=6e-08 W=2.995e-06 $X=26170 $Y=8735 $D=2
M965 255 253 vdd vdd p12ll L=3e-07 W=1.2e-07 $X=26175 $Y=23260 $D=2
M966 vdd 250 220 vdd p12ll L=6e-08 W=1e-06 $X=26235 $Y=16170 $D=2
M967 255 120 256 vdd p12ll L=6e-08 W=5e-07 $X=26245 $Y=22145 $D=2
M968 vdd 254 256 vdd p12ll L=6e-08 W=1e-06 $X=26375 $Y=18030 $D=2
M969 vdd 255 253 vdd p12ll L=6e-08 W=4e-07 $X=26375 $Y=24100 $D=2
M970 180 255 YX[5] vdd p12ll L=6e-08 W=1.25e-06 $X=26375 $Y=27295 $D=2
M971 vdd 253 YX[5] vdd p12ll L=6e-08 W=1.25e-06 $X=26375 $Y=30855 $D=2
M972 254 220 vdd vdd p12ll L=6e-08 W=1e-06 $X=26525 $Y=16170 $D=2
M973 256 120 255 vdd p12ll L=6e-08 W=5e-07 $X=26525 $Y=22145 $D=2
M974 256 213 vdd vdd p12ll L=6e-08 W=1e-06 $X=26665 $Y=18030 $D=2
M975 253 255 vdd vdd p12ll L=6e-08 W=4e-07 $X=26665 $Y=24100 $D=2
M976 YX[5] 255 180 vdd p12ll L=6e-08 W=1.25e-06 $X=26665 $Y=27295 $D=2
M977 YX[5] 253 vdd vdd p12ll L=6e-08 W=1.25e-06 $X=26665 $Y=30855 $D=2
M978 255 120 256 vdd p12ll L=6e-08 W=5e-07 $X=26795 $Y=22145 $D=2
M979 vdd 220 254 vdd p12ll L=6e-08 W=1e-06 $X=26815 $Y=16170 $D=2
M980 vdd 257 258 vdd p12ll L=6e-08 W=1e-06 $X=26930 $Y=8665 $D=2
M981 257 258 vdd vdd p12ll L=3e-07 W=1.2e-07 $X=26940 $Y=10635 $D=2
M982 vdd 255 253 vdd p12ll L=6e-08 W=4e-07 $X=26955 $Y=24100 $D=2
M983 180 255 YX[5] vdd p12ll L=6e-08 W=1.25e-06 $X=26955 $Y=27295 $D=2
M984 vdd 253 YX[5] vdd p12ll L=6e-08 W=1.25e-06 $X=26955 $Y=30855 $D=2
.ENDS
***************************************
.SUBCKT RAS1024X16 VSS VDD D[1] Q[1] BWEN[1] BWEN[0] Q[0] D[0] D[3] Q[3] BWEN[3] BWEN[2] Q[2] D[2] D[5] Q[5] BWEN[5] BWEN[4] Q[4] D[4]
+ D[7] Q[7] BWEN[7] BWEN[6] Q[6] D[6] D[8] Q[8] BWEN[8] BWEN[9] Q[9] D[9] D[10] Q[10] BWEN[10] BWEN[11] Q[11] D[11] D[12] Q[12]
+ BWEN[12] BWEN[13] Q[13] D[13] D[14] Q[14] BWEN[14] BWEN[15] Q[15] D[15] A[8] A[9] A[6] A[7] A[3] A[4] A[5] CEN CLK A[2]
+ A[0] A[1] WEN
** N=414 EP=63 IP=2298 FDC=118037
X3 VSS VDD 4 399 405 411 65smic_062swl_svt_edge_v0p0 $T=109215 6555 1 0 $X=109090 $Y=5999
X4 VSS VDD 5 400 406 412 65smic_062swl_svt_edge_v0p0 $T=109215 22555 0 0 $X=109090 $Y=22370
X5 VSS VDD 1 403 401 413 65smic_062swl_svt_edge_v0p0 $T=110455 23755 0 180 $X=109090 $Y=23199
X6 VSS VDD 1 404 402 414 65smic_062swl_svt_edge_v0p0 $T=110455 40755 1 180 $X=109090 $Y=40570
X7 VSS VDD 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55
+ 56 57 58 59 60 61 62 63 64 65 66 67 68 69 36 37 VSS 6 7 8
+ 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28
+ 29 30 31 32 33 34 35
+ bitcell64_dummy_620_VHSSP $T=1365 41705 0 180 $X=0 $Y=5320
X8 VSS VDD 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 101 102 70 71 72 73
+ 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93
+ 94 95 96 97 98 99 100
+ bitcell64_dummy_620_VHSSP $T=1365 75080 1 180 $X=0 $Y=74795
X9 VSS VDD 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55
+ 56 57 58 59 60 61 62 63 64 65 66 67 68 69 36 37 VSS 6 7 8
+ 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28
+ 29 30 31 32 33 34 35
+ bitcell64_dummy_620_VHSSP $T=80725 41705 1 0 $X=80600 $Y=5320
X10 VSS VDD 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 101 102 70 71 72 73
+ 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93
+ 94 95 96 97 98 99 100
+ bitcell64_dummy_620_VHSSP $T=80725 75080 0 0 $X=80600 $Y=74795
X11 VSS VDD 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185
+ 186 187 188 189 190 191 192 193 194 195 196 197 198 199 166 167 135 136 137 138
+ 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158
+ 159 160 161 162 163 164 165
+ bitcell64_dummy_620_VHSSP $T=110455 75080 1 180 $X=109090 $Y=74795
X12 VSS VDD 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249
+ 250 251 252 253 254 255 256 257 258 259 260 261 262 263 230 231 VSS 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229
+ bitcell64_dummy_620_VHSSP $T=189815 41705 1 0 $X=189690 $Y=5320
X13 VSS VDD 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185
+ 186 187 188 189 190 191 192 193 194 195 196 197 198 199 166 167 135 136 137 138
+ 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158
+ 159 160 161 162 163 164 165
+ bitcell64_dummy_620_VHSSP $T=189815 75080 0 0 $X=189690 $Y=74795
X18 VSS VDD 69 68 67 66 65 64 63 62 61 60 59 58 57 56 55 54 53 52
+ 51 50 49 48 47 46 45 44 43 42 41 40 39 38 37 36 35 34 33 32
+ 31 30 29 28 27 26 25 24 23 22 21 20 19 18 17 16 15 14 13 12
+ 11 10 9 8 7 6 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 D[1] Q[1] BWEN[1] D[0] Q[0] BWEN[0] 352 351 353
+ 354 355 356 357 358 359 360 361 362 363 364 365
+ Y8_X128_D2_BW_620_VHSSP $T=21205 0 1 180 $X=45 $Y=0
X19 VSS VDD 69 68 67 66 65 64 63 62 61 60 59 58 57 56 55 54 53 52
+ 51 50 49 48 47 46 45 44 43 42 41 40 39 38 37 36 35 34 33 32
+ 31 30 29 28 27 26 25 24 23 22 21 20 19 18 17 16 15 14 13 12
+ 11 10 9 8 7 6 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 D[3] Q[3] BWEN[3] D[2] Q[2] BWEN[2] 352 351 353
+ 354 355 356 357 358 359 360 361 362 363 364 365
+ Y8_X128_D2_BW_620_VHSSP $T=41045 0 1 180 $X=19885 $Y=0
X20 VSS VDD 69 68 67 66 65 64 63 62 61 60 59 58 57 56 55 54 53 52
+ 51 50 49 48 47 46 45 44 43 42 41 40 39 38 37 36 35 34 33 32
+ 31 30 29 28 27 26 25 24 23 22 21 20 19 18 17 16 15 14 13 12
+ 11 10 9 8 7 6 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 D[5] Q[5] BWEN[5] D[4] Q[4] BWEN[4] 352 351 353
+ 354 355 356 357 358 359 360 361 362 363 364 365
+ Y8_X128_D2_BW_620_VHSSP $T=60885 0 1 180 $X=39725 $Y=0
X21 VSS VDD 69 68 67 66 65 64 63 62 61 60 59 58 57 56 55 54 53 52
+ 51 50 49 48 47 46 45 44 43 42 41 40 39 38 37 36 35 34 33 32
+ 31 30 29 28 27 26 25 24 23 22 21 20 19 18 17 16 15 14 13 12
+ 11 10 9 8 7 6 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 D[7] Q[7] BWEN[7] D[6] Q[6] BWEN[6] 352 351 353
+ 354 355 356 357 358 359 360 361 362 363 364 365
+ Y8_X128_D2_BW_620_VHSSP $T=80725 0 1 180 $X=59565 $Y=0
X22 VSS VDD 263 262 261 260 259 258 257 256 255 254 253 252 251 250 249 248 247 246
+ 245 244 243 242 241 240 239 238 237 236 235 234 233 232 231 230 229 228 227 226
+ 225 224 223 222 221 220 219 218 217 216 215 214 213 212 211 210 209 208 207 206
+ 205 204 203 202 201 200 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188
+ 189 190 191 192 193 194 195 196 197 198 199 D[8] Q[8] BWEN[8] D[9] Q[9] BWEN[9] 352 351 353
+ 354 355 356 357 358 359 360 361 362 363 364 365
+ Y8_X128_D2_BW_620_VHSSP $T=110455 0 0 0 $X=109135 $Y=0
X23 VSS VDD 263 262 261 260 259 258 257 256 255 254 253 252 251 250 249 248 247 246
+ 245 244 243 242 241 240 239 238 237 236 235 234 233 232 231 230 229 228 227 226
+ 225 224 223 222 221 220 219 218 217 216 215 214 213 212 211 210 209 208 207 206
+ 205 204 203 202 201 200 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188
+ 189 190 191 192 193 194 195 196 197 198 199 D[10] Q[10] BWEN[10] D[11] Q[11] BWEN[11] 352 351 353
+ 354 355 356 357 358 359 360 361 362 363 364 365
+ Y8_X128_D2_BW_620_VHSSP $T=130295 0 0 0 $X=128975 $Y=0
X24 VSS VDD 263 262 261 260 259 258 257 256 255 254 253 252 251 250 249 248 247 246
+ 245 244 243 242 241 240 239 238 237 236 235 234 233 232 231 230 229 228 227 226
+ 225 224 223 222 221 220 219 218 217 216 215 214 213 212 211 210 209 208 207 206
+ 205 204 203 202 201 200 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188
+ 189 190 191 192 193 194 195 196 197 198 199 D[12] Q[12] BWEN[12] D[13] Q[13] BWEN[13] 352 351 353
+ 354 355 356 357 358 359 360 361 362 363 364 365
+ Y8_X128_D2_BW_620_VHSSP $T=150135 0 0 0 $X=148815 $Y=0
X25 VSS VDD 263 262 261 260 259 258 257 256 255 254 253 252 251 250 249 248 247 246
+ 245 244 243 242 241 240 239 238 237 236 235 234 233 232 231 230 229 228 227 226
+ 225 224 223 222 221 220 219 218 217 216 215 214 213 212 211 210 209 208 207 206
+ 205 204 203 202 201 200 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188
+ 189 190 191 192 193 194 195 196 197 198 199 D[14] Q[14] BWEN[14] D[15] Q[15] BWEN[15] 352 351 353
+ 354 355 356 357 358 359 360 361 362 363 364 365
+ Y8_X128_D2_BW_620_VHSSP $T=169975 0 0 0 $X=168655 $Y=0
X26 VSS VSS VDD 1 VSS bitcell_dummy_left_2A_st_620_VHSSP $T=110455 40755 0 180 $X=109090 $Y=39570
X27 VSS 224 225 226 227 VDD 1 228 229 230 231 ICV_8 $T=110455 24755 0 180 $X=109090 $Y=23570
X28 VSS 216 217 218 219 VDD 1 220 221 222 223 ICV_8 $T=110455 28755 0 180 $X=109090 $Y=27570
X29 VSS 208 209 210 211 VDD 1 212 213 214 215 ICV_8 $T=110455 32755 0 180 $X=109090 $Y=31570
X30 VSS 200 201 202 203 VDD 1 204 205 206 207 ICV_8 $T=110455 36755 0 180 $X=109090 $Y=35570
X31 VSS 256 257 258 259 312 VDD 260 261 262 263 4 1 ICV_10 $T=110455 7555 0 180 $X=109090 $Y=6370
X32 VSS 248 249 250 251 313 VDD 252 253 254 255 312 1 ICV_10 $T=110455 11555 0 180 $X=109090 $Y=10370
X33 VSS 240 241 242 243 314 VDD 244 245 246 247 313 1 ICV_10 $T=110455 15555 0 180 $X=109090 $Y=14370
X34 VSS 232 233 234 235 5 VDD 236 237 238 239 314 1 ICV_10 $T=110455 19555 0 180 $X=109090 $Y=18370
X36 335 336 337 338 339 340 VDD VSS 329 330 331 332 342 343 344 345 6 7 8 9
+ 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29
+ 30 31 32 33 34 35 36 37 200 201 202 203 204 205 206 207 208 209 210 211
+ 212 213 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231
+ 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57
+ 58 59 60 61 62 63 64 65 66 67 68 69 232 233 234 235 236 237 238 239
+ 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259
+ 260 261 262 263
+ XDEC64_VHSSP $T=81965 40355 1 0 $X=80565 $Y=5605
X37 348 349 337 338 339 340 VDD VSS 329 330 331 332 342 343 344 345 71 72 73 74
+ 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94
+ 95 96 97 98 99 100 101 102 136 137 138 139 140 141 142 143 144 145 146 147
+ 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 168 169 170 171 172 173 174 175
+ 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195
+ 196 197 198 199
+ XDEC64_VHSSP $T=81965 76430 0 0 $X=80565 $Y=76080
X38 VSS VDD 376 1 377 SOP_DC_X128Y8_620 $T=81965 0 0 0 $X=80565 $Y=0
X39 VDD VSS 376 337 A[8] 338 340 339 A[9] A[6] 349 336 348 335 A[7] 329 361 360 330 A[5]
+ A[3] CEN 331 CLK 332 377 1 345 342 343 344 A[4] 357 354 70 358 WEN 351 352 365
+ 356 A[2] 355 362 A[0] 363 353 A[1] 359 135 364
+ Logic_leafcell_X128Y8_VHS $T=81965 41705 0 0 $X=80050 $Y=39290
.ENDS
***************************************
